//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
SV1ZVBBiX/9se9hQ37sGNGjTu0vl/z8t+YE5uhlWKtxwbPZCzn7v1Ji0c9Em2E4V
fFor4NpyWcW023wyBRuZxTsFATOeuRs6vJjaRa0NRUI7tY9zirUQtvp5/FF7ed7q
h9ITgUuQP/sgbiu6YgjWiLz522tDo3gYtz1kZV52U7JHOvsFWyYaHlF0La5hKV8q
MyeZyJcXiCWRpEm3qHDdis7wbiChtFPSO0+nWT98wvaJIOdwPKv2XT9brf4GVh3L
yWNQTKqEtT8DDqzXBv2ytta9S2dKm+AtC3BivUS8BVE2qghNp7lK/F3DbWZNd9UF
2ZhvMf7FKCUddSVp5GlGhQ==
//pragma protect end_key_block
//pragma protect digest_block
3duzmGwHUOX9V/HDF6Q8ctgf3Bk=
//pragma protect end_digest_block
//pragma protect data_block
BaWnQZitA2wGmlNHJzRAt1fDih/eXv4pNdnquCSw+Yrzsf8AnYyAz07rwd5M3mqK
nQr8HE5Gb//tyCYva726qovBaTB6RoQL+Vmv1IikwMvwSCZl5fZu1PP0M5csssmY
8HIw26OL+d8x+WS/KjXKGwogaxxLMsDBY6Li4adxX1kcaWQATTLTgvLZhGOYF8ND
5dIAKts7lq3xotCqFDVf1Y+LMo7T/H1LfDohbfV0AiMzhlwaE1qB1jPRsNpdcsGq
JqkZ/c/RuO7F6czPysFg7seK7LAi+dwTYGWDtLDx/RQTAIaYlrofw7ShW59hDL4c
nmbsbNI3Svi60LG4vxDyiw==
//pragma protect end_data_block
//pragma protect digest_block
Z+EblH0fI0P/4xRZX+uhzOmTsto=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
XddCncQ+RcPyG5GK8RLc1Y6wDkmyqelIan1spn2d4zzC4EaZ6HTkJpP81+VVfnw0
7H1VxZoA76JrVsbvok8iNnopuwnDb8Ayh8HuT0z0OlRL7nbYS/1QzATuaA/ITbJV
4VrQmqAVPfQLrpv5pRnCmSdz+2g676a9zGq9We3uh/uZZ9ArbRFpNMBoV/eNQUgX
SXhnhAHewX0CYgF58hxe1L8f1HHhUNd1vozlk4i/EokJ1RjndPgWJpz/zADmjZZL
89aDRHZbJUIuPIydJ/fbcrClS2rtznt66iUGR4g+9ZWKvkUUq5HoXe7ozI9U2+/K
dCc39EnPQ/YIBtfS6AycCw==
//pragma protect end_key_block
//pragma protect digest_block
rX0wr6Jie2lfrBhgJkDqFASagGE=
//pragma protect end_digest_block
//pragma protect data_block
sQ1O0sVPI3bbNR2iYLqpq5YY0GBW55y69YSAEt+SfTHWbzDNl8WgxYP5YWua1B7g
vWYDnF8d7fP9up66tBQTTtcsSm2XqbJrtL0CftBjVPy9xPhho21s+DuRHRURrfRq
lYbBdujdyBKuGTLyn81+C3Tw8pYGfizPBQMNY8icj8rUaWFyKOk+aQXCvX+QK+UQ
Q0h73JHKeAVqrw0PPA1FuCHO7tMmnctSY64fxDNJ4os0MEOUQI5HmIoDSccuCJ7v
HKtqPDSVY02w5qJdvutdeRs+tnU1rDB6cKaMVPrTNdqr26gmcralSf4+Fpz3hKoE
LQZ4qd1PBIlABEyhaT6jWA==
//pragma protect end_data_block
//pragma protect digest_block
DMZwznlngX48q5cW+0b4GLPsc6g=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_FD.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
RXHl2YkcKsp6zs3Aezt26+TRYQX4GdPdtoggnl+1xUc9LmSGV812L+uUCsYB6gnJ
6NvhHX+KE+ppjJRPRn5mwB26MyXJaNLHe/Zf5f2hUoGPq3inzRqi/eGj7QmWU6kk
lmsFc6bEkA5j4CwERLIdWKOvE3xud+baJemLtx0uScyNXgSJLQMI7v6rkUcHpIOK
iKnX2bfbZwx7W8cDpy4JsH8DRGIGw3X4+6ASbFFF6JgAVKyy2hYI5l/U7FiXfnAk
2a2fZHi+jz8qTxH2Nv2vGa3NbvAILIUoplV6NSPWEVtg/0tMnjezcW9hRcJOeQ8k
05NltEkG9115qXiBlVRT6w==
//pragma protect end_key_block
//pragma protect digest_block
ueNqQ8PcOIT7hqFSnveyT/kHPqc=
//pragma protect end_digest_block
//pragma protect data_block
JVDxAx+zkjMCMKd0p2Gy7beKa3m5kZ2JVKcVok8oxMel8aItPkRPIwXDuFV2gESQ
whe8dk11xfbirWeaFNshoc6R0LNxac5af3LoN9YYOp4Uj+H/Up3iGt7TaJOnpEgh
N1YI5YYu57FopLpbTOvahypN0tu2HIGdVCmsKBDfIBlzqdvFL6TwK3DNUilRGaQR
Hg/ZBkQA7xKpOneO0HsAWJK5N4l3qCGNMGYiqjIbrLZhWIAyya0TIfMEqaif3+PG
kAxa/OL27MMnp68hyQgvC4Yh0I7V6nMUGkVW+Gejg6jWEwuPt9tsDWxvoMH9i90b
FQ5y+NZkQTuI2DieRZILGFfM1j7KfadaPdAwr8UDnF+AGOqDYC53VvqsPC3D47cF
UAYoO8KiJRA0EvrhhUwNO3Xz27gYGAJzxSmFaJdOJw0N5hvsL7Npy1f3SY4Wt1+c
E0eVJOK8OHQYg5EC9yRrrYUChMRqNbnvmONFOubrXA6AW/f/JVvHiE9KRyMpNf96
gfXbg9Mvv8qw3Q03jCCEp9iBbWzuBeNKVnuU25DRtvtBZAGO6vIPxUVX2CHSbm0i
rAPof9SCi26/pYnM/vuuWw1rVi6WYLf5a2+7gJMR0dYfX6CH85RScHUcGj/vCFJ+
6AH37C9DpZW83zIlHIvkUr4l+nk/ga2yu5j8A4HMR6f8OYOPoouEB+ybc21M6VQC
z1mURZC02rS0S1NBbiwIyACHCtQPioxFaRMceJ695rA/+Wbj4IU2398tZ62A9bUe
5HzZcA1gY0p8oFclsPyJugy68ZmLIH3gPB6UEQE/SucF4R/MJOyG8hXkDMa4wBCA
DI0SaFmBr4j87Q1k6MY2GpPM2Htk6N+gnF6+k6bquoSXuCbBafO4YejXvWPJbetS
BY8ijiOK4u3WjieY8L6kAisilE3niwdFiBSTLjwhbuSW5BZ3yXUnexsCT/kjd5QK
yDAi2W1pTMzipjqW0VBUCTdhuobv7C2819uQjBNOAiE9pPbdFODeujIkeMJ6jrCt
0rM2FodShkxV6YoU97+L7FTu0OmYFiUkIp/nOM5ESHhC675JpQz+b6Wh7ucyyHYX
BROOp+PM/xBRS+MLjfTHoCzGc5N9EwdTtzRqxfmUSOov9nW9HK/Y+7WUbn+IlkX9
/rWFk396V0nMsWf1SVGY/0gseNoRJt0vYSfvbpb2NR6cNBgwu2vdZ4Z7r22Z4LyW
OMbMdRrlInqn+juqHaK+kDKByktWkcvHcJjfqXOW20eRP63XxHyJVo/QFgb0t4L0
ieUT4BFW8pLLLWiWRaWCV0id1Cr/Ag9d8v8vWMei9ggQ1sCjvbmDP92GEifrFe8C
2/NWR4yRDc2gvWRmXbhya4sM1mX1T25RZ0H7aIJGAGrkf9nPbZWAveFM4QkVoadJ
8bhQJAdns/dIJckKkD4ms+WcJm5rz4NNg28pXtXx1DO/pPZTPcNOILXALJNB+1rz
pfCBlpIhLg2dS0/qd71Je2WWth6dCQ6Zogd/SY3M6TlMEQeWXTfgjIj7ysPdNKjP
KmNLFXuL+SX6/UQWsyQZ4LqEC1HxojyukJXNX+xLeQMUqNZB6B8kRoNPxzRJ4SfI
mYT03EGrC9FqyEZ+5hV5/yKexuZFs0pc0vHX2Gg1SuNpgAwTnX8RYBVeEn2h3yUH
n9LdpVdayi5oYOChRllbFKDJrgLVXJlo060LNW7clJ9o9s4nbZ5HXe3hBS4pJAyZ
a0Tn5G1a06jsj6IqxINocs2Z+NSB0vevRj5FCMWRLtvsO6GyjoF13Ft6JRYIYRkY
satGAEWE8LxPnj9K2Qd2vKg0w0JMQm97NJEavR9+DmoMbEuoecJbuf4QYUeiLqwZ
7QvcmCcg3CRodLtc46hlHXX9GKSgCxJH5n0jKZVEW+HoLhVMeFVuysgesSOBak8j
fYa0aWJ8o2BXFQfsOJVgpaSMTrJwv8+FfxaLd/E/HL5nrJ1jj0nxQU7nKt6ehk9l
UT9gxDct110C8v8N9nFTzfzhBwrlbYxu/6sVP564Gg3NB9hapt55jUvjR6VEGm0w
VsTY+MyRKFFMPmJUz9I51B2qvfR/e9utJ7Fv7xGxhWMn/WtlMTzRfKLujMhLdqxd
zQ+chFfsBzQiK0/VExpGqiGzt041d8VHygbGC/IhMd1k2KrKN/xicyELdHZpKB9p
gb/DslgC4NyXMi+TgsWtOi2B2xopXqqvVNK5gzhZ2Q5TIrUcrR7PzlM5Uai+V3vJ
jOoaUbRkVdirR/gzhl7NCbS8yG7SdVXOLpFebNpMm5CH2TX7CDKO3Cm5+ieVtLEk
ESXTeYON8gm6U0gL3mSfrvt5Y32EHeMbu33ymVBww9RFocaiJmMJw3Ad72eb0Jf0
8AZgunFrxguGV8BhJ6inQNyUcKHLgJjzCeLWShsdlURiX3zRhmcmmVmDN53zN5IA
QjxNhBul65Dmu/CjMEMUTVr/OtxB8MFUbWG2sQQkSRw3+YaPZPaz/zerMUA7jxrP
vjY/NILio9V8/fo/GytINfw3JfKWaY69TjsSmqBAOfeBRhqQbyLLhdZf17iej94g
2i6os1gXAzKGmFy418VdrXCVoYQOLSsO4WMF72111+hd9QE8MezUi6cIbptsPbxl
M1tppUrMb27lwSsPHircZWXUkYF2ANHjhmzdyD1j/CI7EEAk1tttLCtP/5U5wPZX
gFiRGWDPH9JJBtaNx0pmo/7VsmuMQNWdAmuS0vs8RZiJZfcGGwBSXaXLfp49nTAR
kl0wQEsDN7aOogJkOau6pzPiddt528ggNhlSJIKLU+2rUKUeuhsVr7UXfKjUjCSs
/RKwRG5Iba3VL609Bf8MQFiggOhbspzyDY9JuMS/7DZS6KRMxvkC97RnjMjj9xR2
YEN5+dUS6nGyMHffRSpTCzjljMf0wEUDyYKZFDHWDWh8+IgX/wrMYZFQEbOuYSIH
5gyqmeeB9Npw4jndiQsNJSdqZF99WjsQTWksIJwxrwLGhsFKpo6VEsWBX17ZFClF
M1zs26cn/l742zV+t5Ty+w9dG/GxtLLLAQBsfL+M9ynE8gqBfrBpEJSj9cHST9dw
LQe3xRx9UYwA+jroxpqgkST88Y7lMkj3Hny4kOyFaImGrAY5l9FkUtSPMELIpMTS
9RIkZtGSbSo4S0KskJ2KG2iM/sXn8HIugetDrjc8fx/1SC+mOl4T9wdne4X2n2tN
aN22VUMBrsdbwIltkkbkBL93fUhyMTRdYJA3DZ8ZC93n55P+wLdr9Aee/pU22m/y
pcw3DLxN6hdhETY3852jE9gqgFmYo13FVl1YiuPGkU35H+FiwPjL21mzS+1HljTD
MyYsNHKe8S52HjiEg98XKMWRaY309tUkMq0riKDagLl2HcBEqbXgJw1lE/VIhscq
Piy/tzvkyAkZGM4CrNvu0MrFt6Eb0shv0DK6uacua0skJ6IPIRwCAFjnUGWWSgxR
Y/LFdM90OjgrXApXoDFrVjzxMKWaPXb0mJP2a8j2ac73qU+nkUdb8ATcXEwbzaie
jhliQNsJPPGd6wn5YyGdQc6KjwS6r6jYGawW+62GQS42a/AjvRSTXSW/M2at/go2
FwgIL/mFsA1whabACcTAoEMJWw4nbh6uqYTyhCg/fzMCZTizwiNHrBZEGABB+7JB
3Dyk+47CnLDWoaBN3lZBQDvQihFw5+bVcnv5JNbj5+iaTK5+dkjjNh4RWFuP3LOs
kUH8oDHCX7KZEXy1YGVkSpDDKo6CfyxBvRjy28iRP5HDGop6Y44HuCVqtb6KU107
UPvDEl7hlAt+bZfl/qYD+HWUGxuzSUCGxyeT5VwyCDCyvLKLFvHQCSVsoTYGgXgG
jQVtiJeRAB8aXD9dJOFxr7A1cyYsJl3PHESiHiGWnjnci2wDa1Wzugcdu4oICU85
hmu+2gQK/g8qmgJTjc/Gx6wGlIIGLBn1gfprQTJG1rbcSYERtlMvrCYrXsk7X+Y8
aNfnGb9gOZddZoXV1/Ml8jjxE1hT/uYpqtPnCg8mhEpaMWamPLKzFLg4JCKZcAnL
bhXhzgMDUALLIOgTORpHA1xumiz7NF1RETRcu2MWdaf8jX+1nZ6+gLx9c9KCUu8g
ogkFprrCw4hqh+Uc6L1nPpgu+F1AYoxkZUrr7B04wovUQfad3ZhvP1owwiUdhBxM
1rf7EXUcjBYPNqeE8y5QxDu/pBSD+zKSjFKcw6IGH4lpHS4afsmqBIjcpavhklBj
H4ZdCYi+aJvtrc7k+hgJBdXTu6pqU6w6wpUs05Jg+BttAEeLsupLChmZv7MDGd8H
CqrZ2DxK2JuDUejCrt1Uv4q6DvoWnZaVygKGSRTMcK9sd+ijuF/nfJPaLXEmKqjK
TDHeoKrMwKiDsUHT5dJgyzY7MoQ37j1fbzmZGM/Qr/VPP/ASd4hpHxYuhHTqRFXC
+Ltn1cix8MCzL260t1DB7z1qCxKtObXtzfLLAhVtL+PAi4R6f3M7YV+AJoeAv8ta
8pI8QONW/fZgeZ9IKWZc9yYvlTuNcZKKZQW223nmKqugrfdysH1LbjjGwHllMIV/
BIerglFi9AErpzM6ay9FstEWmnQGEQRQFqpx+a8fq8KOOXcwAJpQjvKDQgk8BkES
uSYJtrKRrA5ogZo290eGCslCuauClr4L8QvILpT7euMERWj0VFqgxH1QBxectnSV
JFScdVR62A2Twdl3/Cxw2rsPn2vHWFK8MMBMfjqjyz9dpc/ohkcXzG2ckVpBNwNa
DoaGOZT+IGJRTQxfFngN3quFoYYM+rAx3hFWeylpXJ6xYuTz537sMgujW53FVWHG
EmCBoMIM21FxCXa60P2yjtLuA+2VPwYz4n2YiLTPtzNmvzZ/zCK6q8uHazgusKpM
DO7NenEkRrpyLJdMetQs4ktaYyrJUpKCxVkRL9t7WZVhfHx+zbwNZXpNbRAhkCjR
Xa8eGT8lRjw483BxsWARD83+Toe3AlAdY5v6pWciaCi2BKPhgmSBHhmmZju3/+tX
gn27jkGLOk1w3/bIYRDTfcoYLbmLzmG0qDoEdDfm+P+sjGybbQ28pHNi1olTBZOW
C7tY9iRR+6rFs7BWaaVhgBYa5YZNdr8IHGQmHDdWrpX4AHjHOo22pproC0imcpgI
ZAa3M9tmTJ4vpyngCr9gfXds+/ji4TnaCstYy7F4cPvLgfqlYQCC/fyicJZ/PAOf
cIxG+yiYaWwTFJ+l6FgTsQ3WSmAuqoCTuktARjHLH+vVdiKKgFg2MH5JREKWQ2y+
qKGb8Wzolv6J+JKwIZ7Xsr6FlA5nYiwTym970aq4YBhjqpEzLmyUkGjGH59+LeVW
2AfpCvlbNvutlxN2ezlVQKNiKyEpXw+R1R9HFte92U2byLxySnspo2NKUuS0DgUW
aMDrJ8JxBZVj5APQLRdVHXEe8c5ra40NxbKe+lNZajshzNBkx/0IpOBrJ9fIdJyF
a5Dg5HgVf2kdeat2vWG/s0zP7cR9QKd+JpeFrG8fSSj+GbyKyHEI3ZLHeVM3Wyu/
TPWOgJmrvHZCme9fampuMMhpGgYHI8Br3Gz/QhG1NU98SsYf5tqhLRZdRw/N4fWo
3M2smfpE5tOEATSjn3sFLcl41BzDv5yWcmMR5ubMailMq77d0bJv/Erio3POcDLM
fEqd9v0l1nxrWtRNeDesuFrSN5zD9uPk7BTjJ0jfGcoQ8dFSC/VN+HTeqepAvLnU
4BtoAcj0vCVgc4b5kQXdCRugbuyXCFSJYaWviuhkAVNsmypnm3cDRfE6DeAUTjTH
8Xs5gzuUwqvSoTKFDEnICftYgZtSUwlVmjAjmxjLkHayuqQ9tR3f2vXnH69B0xBH
ZddiOwTS6js7cH7VszvOZqkIOWPxxqeCMA2AoKn5N6ab4LLoZ4SfNGDHtGa/kmwo
NPPQNizcPfxmCYf7Xk6yvk1N8IWm5VPT0Pv9wNl92cEzvm0wO8+ZvgAO+E5mFmCv
lG8wXdGarAkZchuj+b4EF1s23iv35HHHgqTX5CmwNwE1gU+pAzT71pPAumYeh0hy
fPddOul/bgbyhooLXrjpG3RjDGfL0lDBXD2HNpW+5K+UAVvmbeDg7c+uFmcd67+e
k1ValF5urhm86ERz/lMkL3YyblpfnJlPkvZKZ1LDrshTZtlDoaRNacedcLtQKnZH
MvnkolIo5JsfXH9M+026YlhzgrxNGWaMq2oGOq7BvOtyOTRESFtPRnIo5C61RtzV
cl0dxrFXSvOjTWReS7mSIXDBxQisQP53FVaajQ1s7D1ZmxcJPhS8/5c0+89TOaDY
+e/dL25ZvFtX+b0zjVnEjlIrwzXYWYAhCQaZ09n2AHb9S+NT2v4bZ4rSFLmvTN56
Pts748GcXlW5CR6XvxzEbg6M0B41JvLud3bG27topN2/g8rKgKG6r2aTMvGKDOF6
hbbwUQcum+nm8GU3xnCdRmyM8vBO6aR43fVYeP+SIfIz8sYpa77lWTg5eEVl1BGY
VmvKPeOAnBfizzWEPzSpDrMMjyeqtzj7Kkt2++ByCvoIz3ga8T/FXx0Zn11NrnFT
8OeXRwdyFU6LlIQ9tNZpbVRsvnTSx2nhtlnk//Hm2tEgN+gYeeETkItaJ8Va7Z/u
F+x5VgwzYX8lY7yK35WvIDuKiRuD1Ekv0+ommFdm2pWfNFYGh3wW+yBOnFDGhwWm
HZd/L6pFMXcL1fvSKgvX9UMusR/8JukT0ncK4gN7y22qIPXTVd7pT+rVRDN1vLly
bwrGR8wbR4lGXC4Biex6054rsbXDceAe8eQUjzyXeMcmGzYISRgNG7KsCGBNSP6u
aPgNNQR+vfAxco1pWlaxKOXithWI0wurV2s78MM9DhjulL+ZsagBcRXGBGSbeGZP
cLKT1ZLUu57RZXz/CckoKPxEXSSuRxTg5Q/mojzf/oT71uBZ9OKXbZkt2Yo/8CyQ
iFXxn7/FF4sIk/OVHaetRAKJaZAr6qwjEBbZhSKmWvCFOLGy26RMEj1q8t2rI3Z+
8JIqPx4Ea22aoAmqImW8h+N+qDVZY796Fc5vL0MmR+/PXfVNHAxDnQT8kNC1QUbZ
hg6EUGlVnyKPtO/dvnBtMGq52BY91c1KVlmdBlHdOxXVDsaVxtP6uqlsq75HRmg8
ff/HotsCW016p6aeADrhYwwmg7th7d3H9fqrrDCQwOtcltAyVvmZfcbFL0mD6lUf
EeLZAiG8hStBtd8mjQ0thDuyxXVbccBbcLSj4ORbKZ1Y63JCD+B6N/qQruVUn6UT
lxacdhRb40nKurDagLImSa8OvlBJqPuPRZ9gST9sqkzYhglQNPqYA9KtedIHMjuV
cqHC7sMy/Sj9S4jYlcI6VHm+Y83OPjyaEJ4MxgJQSvlzB02QJq+iY5nehifQHF6Y
Y/ZAFVncj96FJUzWm6UrSRO8PeYIRfIuWgkDKfBLP4E1V2077ysWnODSChXjobwU
pQ0v83Ynrw2YVHQvBAAi2GrH2sdK8fOh8/VZlF/UB3LVg4eH4JSOaCwYfnbZ5jhr
PUlj2OqLHGO1O4dq/FL4bKxy0bMxExVF0tymnfEekocza9N77tn0JMfQguiEXj4i
rMzs+hD8EuhO4bL7Pdb24ECvI4IXnFaYSEymZ20+qDwHylbay/gVfC3dukBeqyJq
UJWdTKdTzYf5aw1W8DljiTZvEs7JwTrRjWAKX9VFQ/12DdNG+mUovKIUSb6oFqa9
bec7wFsHJSEVuvZ0z1Af3rzlS0GgsW1Ar930dUWe4VNYf2zoAwWhERDaF1oUgBdE
56z+5mNnGPhNZLY2J6cD8bads7AFeSHsggXI9XnoyV8433SA14nKQIaMPlcvOH6n
dI00x6/ghLhD5zYSyyTwM/05H2CPjbVCWN9UFvEy+OfgBvYRD38ZbKnVuKpgvnbT
vGD+ZESIdh40tA1cQBpKZWliJD0gtIJhY6KHspK1ytoIkXKDvbWmRpl2Axx3ue3d
LBYD05LY1nvua3hELlYqz4q+oRI18LO4TKBSjaKWOSxtyg84AHJZX23OD723QctR
791/P/OIfg5duqg0I9qBn6eB/MiLluQqhXo3tTAs+QdbnuR84PpHJhGn+i4sV34T
KqAiYers4Mjg9r+DjQayw7crd5g2khLEMCe1jao455t4hRGCInBtg44TRvxvvmFm
hkvXJuTAihYzYVAsE9glo5u/FLFkl3m1gNXpfY9rZaKFrA7/mPApkpw60dBZ8jh4
NmguoyPFbugZwr/C4YD30zoPBkBRulJYSMGt/ONzbU1/K2/6uxn9nPfJR4wlfU5+
Pomc61CuaWTGYYk9VT3aJMHq+YvVfIv2tyEXf63gLyyOFqNup09MJuRzgdzk6ejW
MthY0scisX6T0KOL+Cz6hk8a59DL58/MQVU5EI2I61KkEPxMrqXYe0YGxdYSal0k
2Kh9lP6HH611iWbmFqdgtLOmVok+kgTf67KAN4Xpe3+3t/F+/4ePeaFznT2FCGsL
a7dNhFcjV0IdwVCuz+fB+EIUhT/pr+ni6+3E1Xz4qV39rx0ArM+AUsxWPjPH0Zki
Q8fGRA0bmBzDPAXcGbEz4/gTeSFTMyhpOW3jyU+H8BhQD2SM2zwFyDKVvoAEvVCU
rXQNlMvjiYooGUsJ+GLDoCFz06D0ozp1hqCZaPfIYhpcfbv8iRZvxjkCB+b4Kg7N
uUpjEQEzV/aNyvpLLlfDih9Zhz2sJE+2ilRD1TeklgQZ2Oao5DxK0VT2K5rMAxeL
ivPD4vvTIBVNRAJVyGosaXJ1a/igS0tcbM0u8ObUsZYIz+SnOeDRW+ixFwj46DNd
WBpt8eS7OCwVSWFN5OCO9hUQP+D3v7c6JFIFj7uH2NRR2InOK3OhZ4pf58Brq4m6
dXJrGz4kcFjNaIrLjay/jGAPe6GnsFZggGvahshWFctPMBSYswN7m3cW5ZDjiAaM
d3jrrk67HwYrPm/aTtqEZCdqrQrdvWQ1dLwSN211/mg8aHv1cJ6GAMpHVKWM2iyZ
T5AxzjgCKrBhoeTZ6Wpos3AyrF2Nmy09C+C6LYuEEXjVrx6mLxY1Id0ehNWYlB5K
sUgjzsmJqsiJncjTPod3e2WElj+dIq1/8fbpcvTxN/J9u27tVObT76dkns6AlWYX
yaWPJmwOiLdK8nLI+/4awsKjxNXzBDPXznl0Uh/OAL3GGdmL6hFz6Hsiab/T1jT8
+ETGTxw3w2jbFIx1dJcrje4JE861dFgJmYM+gu+GvQ44mvvI9PfaQtZsBz85u/JS
9ahGbX5CJRRujFgl+cYDvNgVN4ySG2BGqkK/2bUNTAgblNcfNc4JlPni1gyTwrm4
wiXXM8DcJh1FiP3vcfUkSOkLitZwLVYs2PtAVQxkYb8awc3ZKSQKJaqC83Pbh/q9
XViUATahGH54ceNHotGOefgOTvZn3HcXCnKGLqBczxxeVHzhPvEj/tVM8yOqJP0F
C5h2jNUgmR29L8JbwvWp9/gRvuePEB5nEx6CJlShpAQloY08TMl2tCbasiLo11uG
e4jGAYvNoMmRGTcm5ReIRxSSMAwxGr92neZMGWHFR8QiLdaIdmy8ubsu01ZI+1v7
d7FoJYsDiCaHbYRur6YWaske0lGTRNKzX1lwkLK+k6inJurqKHiwAw7hZncN8yiJ
AoThFL598QToqVRCwqQ1QSN/hrlquAUjFdwDD31dg+WuwB3ZxJD1saUe4jY1qIe8
+MGDljuUKLLBRy8YsYkwHdMRzUztSirRGVsGI0RKNEz+B7L+/rAknvobYlk2A9VP
AeaYHPvpyDx0DeeWcr+WYnDlv/+kqxkS7Ve6yDRrQKWu2FgB8bVdsvD7ME5JlOyg
NbbnLA4UbWJf1ONa21xammaTCYMipuKU0B+3Oo9YOY9pYBh13tdiZrKO0oH3SqB8
WqZsPMwrzEi9PSfGJt6PCIXkjqv2q3OrG+1pk2BXlGMOlNceZQVRgi6FOUfyiLpv
Tlahq1FUOH2Vwm55CfABgjr/plsTxOYKXfYHrba20cb2HqDthWkBM+Uv8A9tKWhM
842arkcjylrX5NazmMHtk9ZjkJs8IZ7drgbaOnoIOptUsgakCq8ii7p+HpOKdQgb
fJnu7tPhtqOr9TkBbzDnE63EHVj3vjYJSokqwP5BtDk9jFD4StHBpcTbwHP6WMi2
7s9NQmC3xO7FNTGa6OpM6UrodjWdLaecLBXP5myQw6WLagb+X31kdxThhBKVSUMv
7OH/d/13gperzE41ZB8sBLq0Wi7sa0nty2hTO0FgJ5mIPK+Nxa6kAaA3X5shey6O
fyk3/worwSSw6hw5dG2AXrOZNHJd5ZX5TWByQ4NFbx5Yx9pkuNa1ZQQC0U6mXKRC
mT+j0HDBe6OY12Ij6/trqhIAEmksu56HTtOTyS1dNh/2Qen3ICtPMc0UKnlonT68
ZbgAPuw/PMqFiLbozw+FzhkQMd+9nc3BAhHmGaBQc/OX/KweBnBYoqX5CybA7usu
58xxCg97+bPrD5wQFfFntvEVWPSLrcVx6BBFp96/HtjCsjhdxTeLi6od9q9tl/Nl
VVFvgTrHrEMbkTPgxH8ZXtvxGjV2xLDWOnCKd2JmLwo7cYPkZrHoEGPjIxuRdH0z
CatKk0gLDdT3MHB7gSOaMkFkLRQuFOq2RBxHp6sdrGd5ly/cBk98VLhzCM+j2IXX
xxgEj8E7GuS+y9o3dhbzkg5GISE3CY8rGf1cHHwwoF7TU/NnANIyCObENuImbZub
DS0PESCixHLdrsG6T4+WUeNF9Agfs9qAHEVHO4EIBhDKzlHd+NUXO5lMj5nuDM3r
0oIuFS6jGw/4rfpi2wzU8TZpIGl3qdMAD3O8aJqmi88JoJOsqkHUs+vItiEX2Sxf
kvp7c+RxO/L/to7ovixaKI8MX0xyZ+VGEGCSLWpIeyINnm8o02/vVSGYF0rYRr7+
qUQlEBOQOnbTe7/jKCQQ8qE5o/W8gh5iZgBJXUjIjVupDyGBKvUYV+bEIasZzT/7
WIZEofW4GE9AHmyrgJwsyKmRt4Jo2m7VW+rgP7QwE+Y9jKoKO443R/UH+tLBqihw
ElwBhtmC/6XNzL5EYY97EnKgGhwcl/PJTuYN1SKq0uNsMAr2SZuzsM0R/z6Ma7fp
6pmZoG85HEPz/wv+ubTjvDUGYZT/WdyR8Rc6TV2LOAEviYNtUtX/kAj1f5kwVBma
Sn8nbVdMosmJws0im+OM54yQIbPNxwNBRNwGRwPLKuJ9cG3v9sTsMP7XVuL06GZ5
Yd8RL+mcEJAHZ3fY570NuZURxgxlJu0YGJf7ql9+gG832kwCBgzzwkoQc2qgwt1Y
oWI/AV+vnS5QSOc2D/SdL0Z++9/VltKHZKgNoLY1Chy166mtYMNOd+M3z2qpqupu
ynKGxQEoVdhDUTgvYRV0wIVMS5nAZO1Q0Cq3rwKN6qrdQvEwLlMWB2OGA227iUMt
KTuLiGjCbGhvZXEKv8+2LH1o3L5FUvM8m1CaFDGdJkGXAB4FnyNqkoG0YrnPd1K0
dl0CDZhpi60ixjglRmSmOBT046yMhwLbA7/ddRuaaSGYDLr6JZDEWzS/YHcES72P
daB+j+/387S4OJPnSfQvMOtB4E/e2hFf9wexV71YAQcdlaIj7WroVSnh/0yiHc7M
758tFFS03Sa5vgtIz+ZBt7dzYTzYUOlODRCie+iFaIawwn3ebBx44tIfa/5UFSeC
zFa9+CwA75E0zBAdmwLUQIfZ1gZ6ObRAwe+J3fRQ1V2yF9ba8FNs/8HlxDPlTXTS
4oYRICB/m/vGG+CxUhApH0+2ip/NDucYXI+f71xQWPlZfDlhtXtDT7GMcXzOIubn
3Xje+bpvTGQvBOYPJgG5IMcyvQKfQdWy27WIAZ6XVqqNis38ABJSnRaWM++EDS1w
AUe7y82W6CXgvLWigZ35DIGBiVi+B0Bj/bgvE3UnuRSTGwQmihS82GgOaprKacEw
R6c01LUUNDcV8n+j9kSAUGPsgXbS+0UPj39iXISm89mLtfBbuzMdZaREFUmGUax3
LY3cSNDsLwm/T6vRhCT1kv5f35/du2UziJ7714Qa3n1nyA7+3AaTaWMOZasakT+5
aFmwzhiJy+w2PgTCksAIES5u+/iZve8x4OLrOle0sH2QC83OiTip8sMLu1KjuLce
DhcupNjethGzo3SdvhgkE1TLUVLj44cNEFq3fBUnbyGt5KHPcmmTV7YUD/nhGz1h
UhI58cMVSPwF1fGilGS/pX8qaFqmHO9ZBkvVHYkrS2ICfebwQu58SR68xTKUQqx5
b2R5MQIv7mYEdoADQDTrE9Iivv+9OjT0WvjwGnzJxwIREAqnz2uhFT5Nz1bHTzJ4
4JUVAhSLkoEh46NH9OjOl0fBdmGPrJA4bzZGFkc9S+RfjpVD++QN/JUXd983Wyw2
EdtdVk6OsTxxGLRvrWJh01dmI7CC1L7XsbYKDFhGBNh/Dr04vX6J25FJzOtr417l
5WHVJuqBTSRtba8UDMR+EGA+HG3BI/N1V243KNLOG0FQIltW8zs9sROKMJa1glHH
+hrOgLJrjhJ1s5pBXgsNP8UEWjsPcb6Dr+iw/v19Bs47d0sn+CSm8pRr/1uP9t8n
RS6bZraHAlYu2xBqkNesRksCXGQYnDXjpCILVN7OrDv3SgSjg0AtZIh6lX76UtKt
fgqY9DG03f0SvZh4kPw+8WagExI757SCw+e+sq4L3LtpJIle9hH3YWfWUNFwLVjG
MWtNxJSUqNJjrwx3vw/cf/wuSpbuO3N+ANfh3lo87SK7MBpnL9b87V5wNcC6Z/Cv
Q6bLCgecrkgHwOQcUg5bP6gFZUZ0OuQvxwf24LW1pRMJyIE0+tKtyqyYWtgJFF+q
aGrsNUgSIm9vqv+Qt85HqXQwZR+QJsz4c7XC3JyPYYCnjKsEf7YsAS3iNjhuRM99
iSzVzqgncjK9LW2DHnM+gGqXgcUglQErKed63+OUO9D771kboJb7UOeMD/lwU+4P
16ACCd3hg8RxveC1ta58bsZFA+BlzJa0EAGyQnwcD0cs2VGpe+UG8KXEJvUbrREe
kHSHk8W2vBkZ7QLrhA8YeLQJcUctN4IhxOJsSLAhLnlL/HIhb8qM8/tCYbjQipmu
wRHpn8pR6x2jWhfXx4Q8P94GE6S60mWFzlBf2WczCVrDPeyS0xSA7WLhozsQr3/k
cqIPoWNU0BUd/syj/HJ/VO/zxQ7i9mdKvWwe+XSKZHbgBgO3ahgr15zC9Rz1dU6W
xR5cmYT9iGl81oaHlCcds7EmhJozmMwtLeyvqJ8GYbjS9umVjJCJ58IuhBNom9e2
ZzsuGeCVxYmKcAtLHq8uA4aswcZhnP7bmhvSfKMH2cb22X3p+DbBtyS+BL/FbZOV
FKxVPIg84ii10OVLisjTQX2Wpgq9tDKJWO8ZBBpn3PItfzPkPDS+A5pBMjd0Y6M6
0VP1OD38izhxWjTAYIPW44HZiMAAczRyMMchcsA/XM7lCoDil5oNR+ktzfiT3Oz4
EX5H7egGJWmiHmgUPO9ds+ATd7FICCgS33x+3zK8Nq2SQbsAhcZJZeYUkOBJwr2Y
2osdrwpDpcPMFqCtF9Pu577+e44jlP2dHmMfSiwa3/ijFAgp2H/lAxxdwlqAjZiO
JfzGpwHlF6qxQiXpqq9F+vgmrGXCOmvmNjPwt4v+v395ws7XnH9Cb83sXOxADxum
N2REuKj4gAvaLvxc3iMvKQRzMlWfpetHzIGq5dSdx5zur4SjnN1flvt7/1CCNNkB
EcRmRVEStGlM+F70e9tn/USoUKgsduMQe0LJIPNQXjgkNSCeABiaPTTEDGKzXhaV
o+mnaVxnx3qjBhHJhXQnxKjnJfy4ATQdrXPMtNrdHEYCe2wMuiqUUIgsv1vTGMks
rv1wVLleIx8E0qPDnRRie2Yv/Ro4EWXryRvJHxPtfsR6tzdxQerAovOVEzxtlNc7
mEp5teFZxhFBgFh32klKUA/moP20SOHFhyApvmufX2gNdVaqez1w/Qyo+K3IIFiT
tLc6NqccDZCqK+/WRyJ+K504zx0p3GHhRJS4y0bE4OSrIoog+ft+4UVPbM+EtfWG
/wzwYvnfmEgJNQN2pXpQF/HsSBnvq2Et0WbWjf1QrwEA7yDjFErPpkjrWydKKarl
5pnOisGxzpDoJYy4AkTDx/ze/qxVzROZxqBICe6O/44RF4VPy1Uy+2hUuFjurMAp
YprD1Ozy/ISrY9UEjQyN2lmx1qYfZ1qy0129JyHEfqcbWIyWwY5V162qSmAkAbGF
mU7165j8XTrf7YXAMD7f7fcHSreoRr49v1iFCjO5smeve4iPCETY7ZpaE2ielWvj
6HNvyqPOScJefLbwaUWDMo7Kz+MeWYC9ak3v3RdtgtyZD1H01UAHX3nFNU4ccMhs
G2//pcCeP0ocW/KZrNt8iSoeC8x6Q3YIAZByQXNn2+sSRer1Oc3q948esQGVMIDP
RSgD5f5DUzhimHT29sToBYlvuN4edb2YnamU5rV4LePoOuu6c58bNcdHarihZFjy
2ZV7c1tuj9d4wPqriCKI2LzDJEo8Y+jwCtZA8eyl18MIndLhz5o4VwHe0v+BOkGE
t/JOEnd56IImMZpo8IHHy26/CgsdwkLd1XPydwM6b3D+IP2tm5j2i1uauPy3Ekqf
bwLWrB+uQ9I28fDy/wbZKczsRcEJxyo92xJQ0kgflFlFFZ6+FDvoWlty20JrXsJf
0NAeTOi8xV3bF00iyUrrNH1wv14m8Os0dPYBwshLuipEx09UE/1uVcRGlScu5Yml
NQ2e1uvK8xvOtqVB4fmQVHHs3jzb8ibYc0YVjDbw/8uWuTlwW5uvyXKYF8MTX10G
/Beuxq+IYV4oSx1Irob5gD7ise3JfpT4ByJd52/JR3AJOc+QWUAWJdA128Uz6KkG
YAIYtrZGwZimr7ANWcpgmuN1G9qVS9evYVgGZqGQU4TxF08ykIzrJf17bWI92G1o
Si4P8GYuTCoofVGEDE6uvhZzFS0BnKRabrp1MuzBP0nuTUFjTJEMKoSd3eUDGYAn
J/bfyjgM9l0cfI43xxKfJ1zfV/330HQte+DC0earDJDvp6qYwB+6mOwYbZ0j79jK
77gJfHUOVFyCtoePwfBSW5m4onmZ2uxM0lzxn0l1w7SlinD5/Dzi9fFr+mVeJA1f
z81jEqUIxHT+HydpjwpY8uFItZzr2BrlGrdpVF2v7wWfBo2XExldLtCnILGjybA1
JfVOJMTwpdK6/BWTsZxSaTN6HlhBEgpwwAZz4FPku09f/v/10ZhQCYn8uZXy5/t0
P1LRTp5FvtqTFFEjNILRVMOw2DavbqrELhG7M2gcQBv+CphawByGXV7Ehk8e3gGC
HfIvlOY65lZMJLNnoQumxSSOrfiZzfo8Fpmwy0F+lMJN5OG5KdW6PI1AstSyW5Mc
DAygkXG4rRVMO8WofDkl7eNEQg3Zv9GdB1lpRcJ/HrGm9iuQPvkAoFyKdyKi40iO
KUfu/SwVjrM4HCRzULlqmwV1wISg43gtB3wGaYbeARf6nSLew2brQkqOzGCX7B0H
qvdwwrrpfrURH1ak4W5dfVdSaDXEodSDZpDIWaxyGCdJHjN4KwhxkviSrtN1V7qk
IkacOdAD+Gqzh8RR/IyFX13JR4LmRWJVctn/bC3XFaaEA+q/5xJ8mDcNyvs8lk6L
GbvyhT+FGnXxaAn/iNTx+IxutVMdKbe7qIdQXTW7JwdY4W2rMGC4VJQwjN1+84Zh
CLKB2Wk205LPMUNnjp/lm3iBQcD2msE5I28SOzhin8mrMx4Gh5ISCRKd7UQFfbr9
rC5U+iLmfiO90pfddwnJP/iZzOXjsp7zeTJkOOjAu+XiAsUmWXOgaU87LwP1UGLJ
MXVtsPdK86JvxToYGKdnxeYTA6s4NK51K8NmtXYanqk6ZUVf9/Mc9V79sCCgL+xV
B2tqlL8UO0A9NkqgjN6v7xnEoG1MFbIgnN1LAEjq228i4DwBaFe4gUMA9alLTtbD
1hJCebNI5iDtxmJ4To3HZaeKndjvj82x9ySHu09j2qQk9cGLzgTNU57EddLATzSK
h7OiXFfb67pb2sMCn3sUrqdOj8hqexcXfbmfLuiA4a/2dphMgWBrAOb+XWZmTjuR
g6i8j/y/a27AwSUqWVYGuhaetKSM1fYM0+PHZNJcUbtV9IrMnKL1R6QMV3DCtXOL
mbqS/noJf810ZGqhfHSx46tgeqUfCF4Qn8xm9PR6u8iAmD8AkjqCF+tnFYKke98H
K+4OoEIvHHjgCiFR4VvbWoKifSHc5SH3zRYQaaIat/UuW5onYRCRrDo+jTM3cQOB
MEjRwI5uLooQtfuM5T0cUv2EAj8ny4AMzrbz2Uq3GcdgFqeZInK8mTZo8JvULo8p
HsSuysno47XClaNJOyYVNF3behUrtacMDv8E212oIXHFDyjYtkZziMXbEL5EpsWB
fK3HyUbuZn0O85mvjloh//V8qr0QF5HW/UYsJp980KK0IGRH9mf0DA1FdzN6CdlA
yTTOI2hMeaeAcWqhTpu40Z2Ir30TFeTRB4Yw1RNQcE2Aja4ppuX50BFle6ZZZZRO
/cL5/wOiKuIbmbPiwQsKogygCDBCLyZZ9R7IdktA4DI5Y/3OjwLLtA06GUspqpXz
5b27ybYzJwq5hYfEzcQR85GAzKSyiXs4B/Swq0nlLINPUku1XeuG057uUu/3z/5j
q4IEKkqhQOX4Jcne/iTYUGOKIY+cngsgMUwuMEWm0vi+/dv0iTzslQ359cYD1QFX
lFWDoQ7k3gFKhUaR0f2oZPXF4qvXvr7dql6L63vHmGnU1LcPzqch4qsU6eDJmrAW
bJgfe9Py99fVuXMiI3In8yurO1tTcaWp01rmwZl+t1BIMPgXokvUbZE+/iDOwA+U
SC3zyefi3S3J1j00rj4xqU/NMk0UW2uOvEWj1BSIHJ5bWbCd3yufPwT1xokXHL0c
LIV2w2RIScpVo6VFnWhvr+B9JYACyU8tpy8y+f4rTybn1xaRSoClkF2jvnTd3zal
IZ5F0uoGycH9rJA/G8220YyrExWwtEq14P4RpVAg38QL9ZRrhlzPFkEAISV+XjOP
dPAU4K7Is46bluScRRfDLfln24MkBMBHaeB+zYkJ7Nh9e6+2tF5eOXVzTZsPL794
rVT3C7/tiJVjqJ5kkvNlR1IfXwJDxQgIoG2YA0uxd8Ns1nk51kcOupGScpgkpbVA
p9+5NBfAJsFC3/TitRJvlStdD6AGsfx0wq12poReIUdwo33p1pTvNMzym8o7OZ63
4DqS2YpazFr1afQJ21yqdZs1UwTUcig7PVNqxmPMxiUSd/DdRZ4m2+ETe0vevTRZ
1sCWGTmRJztw1Do1JWrQ9cafw/4wDt9Ck1qFMPIE23S85H+3dhfRMZJHh179wH1Z
VZ7t3V4Yyl3CJqK8bmenUnYk41bmiHHNAGXIzYnF6yPP/i/kkAGGzjNDXaIizwDO
6XH+dYhiv7qL77AXLjoX1XYCA4zcaxHnq9ZlQEK2UG3862GIITsyA5sSmnFVkhPf
VDi2dQEIUv3KFJOC4wZ9fz1DF/in4UQhl2Dj/17+tyCHiTVbGIwzXJd05+j7N7VK
hf2Rxc2ojBVTg3pwud3J/aQtUMexddOkS675E/8s4/pPoqdphTkNvFCtbhsuBxTW
xOYK8lA+8ywuFVkJSDcrdp9jgCzA5MZotanXykbxY258uOvLTHv0TJVIKZN9oz77
hAYRS901NhOQUOOe6HO9sX+ft3732gChCRMrD3lOzkF536o7dvh2cnZWrj7h7dSC
wEnwMFkgCiKZy9ftajAgp02yna9JqTgjNfLTfzyJmnDJiiLyvELfu9XezK2V9ZmC
kCPbC7GObOqA00mod9+ZFq4b2IxH2zXUgljo9V2wPVnNJc+iR3sdbVNHOhNPiqxM
E/PjUk2Gjk8/DJfqUB4R41G+vQUY80QKN9geXYyxg3h9AmKaWQcyvDFAb9jlGwnF
uIkfoLkg5VmAFljMhA9qYWtblcozPDFt1NFZNcxx5+OwBcjkD0CHO6xghoJhIHCI
yoFl2z4tb6rphFXvBpitXdykN5S8rEdnPefngvn5MhZLUHh4bYo4YmcIiF/Xz1xE
woNP3jtU6AwJgASl454ZhXakvUE+sIOJRPouTxtAJ9Knw9rlYJT7KXgpe+0Ls97G
7d1AeuWA89AZBDyxKrvu+mgPt+48d5KplLlCLC1a3Ri7j1V5KSPGwwU5ZaTwFnY3
M/O9AqhyxPHO0bFcFSKh+n4YjHkuUB+x6kV0Z6M40AUXC8ApKsQ2qWozuF01UiNr
RQbZ/ilYfv15ejKj+dnagiXqWS83OMThNdH+4rZb2bF8bK2KpFzw0PGm1Z/2kJj2
WKARN4Rs3sU1CyAC+yA3vHfEsnkNXKKXgFug8ZzKt2T9bXcPNAekW19dx4lgutwo
zsRmSkGTq4lzdFHdAUE7tUCMSDTW8K+BoWcYlDMT9gBcKgCSwea1i5p/uV5zapA6
wiEBalg0YbXhgESp3iZUa7ug3ppeVAP+VWd2xF6HgSQ5CH0ZNtq8yh82/dvRjCno
/Q1Qj7fLiiN2+BKwZsg6ZPIIwg4R8JE6fX7czVMx02cl9/jbplY/Z352Wx5VxZQw
DljxGWsEiWRiF/J89NYfyXW5a3HqaJPy5l8Xrp0MOK8QGLEZjKRSWtxMHecRt2ar
rHsa6PKX39Z38fs7ERLe9er/k2pDD4WsCW83xR7Dj96ZnobBdKz4sBx9OGrga+Pa
pZwQrs8iI33nqD/BOsGoNJNjxQsGGCv2K/uAcjXbHWKmyF4cN5H8bO6VGA3aYCJg
xnUE1iYVeJFlPY22iUVRmU1O/MX9RYTpxeOhzymJCLrvPpVV/Y2PMXxeUWG9ID6/
A1tPiW8buseTc1n1va457Oeso/8TWE+nPn2wx7o8PGgzYE/SQ0WP66sc49yPkgcK
1+M9E0CNfYiH4T30jPwXjhVbBXhyB/KUl//CX5uA++BcO0VG0nj2Qp1kuAzv/tJN
mwK78jVR1LHAwJ1IHAzcIh8nuRkM9Fh+6X1WCGKtuV1QqW0qSwxWv6iS+13x0Npz
3FUibqtAkj1GtAR35wLzof3V118bmtEeYKgCdC0rnbQNieMA/lhCzEaB6gHBdUF0
SgSNVpm+O9EZsK2LzqsByNoU1Dw9ka0CCEg3UUQp7z/CdT47Pyoy+byyeesIp1i2
QqL6McG6zPZRf7XclLn5mOXkFcuaElgW194caRhsmacjaYgnGJp8IAi2dVS1RGoE
NQ5hqfQ5DCEBFM6irVi9aq5WTevSRQSw4z9nuwWfWoiUp3XVImr0tNuJ624i5r5S
JdApiV+y6D4+kFYydjZT6MrhCmRqfweM3n0WbpxF1S0p8jeXIPxQpJ0iNbnGGyDO
5XJ59dLatRLyL+pXRI39isSHN+G+K4SQX+2N0YGDthA7PABnrxw3F1oZn5fzXJG+
mScbOt6/E8R2fZ7j349Kyo1wEt2gUelmmi9HPhn0zq6vvT+jHqC9XE/wBLMlEt5O
QssgNKTqCWsZjqkI3Wv6wIb8piJDVVHyY5bYH58QkruPmgIxkzzZt574Pk6CBTiU
0vSsynDfQCIc+v62bWWc46S1PdUn7B/Qtp9HJAqCS9yuOYcG4WjVfiN7crHFYyym
Yg86N1GELyPbGJfZ5ig7dye4GK3Waz2Qx2bpAZ15HTMDN2a8KnBMFIRoS5W2Wq7d
bD/cQbp8yMsfFzhIYSVUJblnFGDBc/2S9kjvca4A9orOPkLwv2UQIoEtUgdcxtR6
yaFwXa2u6or5o8WbhbPJhQ3d4VUMdfBw6V2ncVx0v2tvEIwMTz6CmGRIfi71e+ne
+I3A5cCxpudYbNYcewjj8bm30v9Q8B1NTlr/TGPyaZ17P6drGCX6B3JxhYj/1o9M
OZPSci5AuwrmZTPz/dZK2jHUu8YJOxCpeoAFOdLsozFREjV/hQ6beRIS4QaxnTzj
Jl2THfPJrhHbytrLZHEFw3FEcfKQhUTgS9KIlzv3T/qFtabZBMxhSJg3cCUSUoGE
f3w2kWO/cQ+/YhMO26u+Z++jjDCCcZFa6so8WAltcDzf3tOPZ5u7IjmQbj4sujA4
R9PW1GPwSXL2ds8r/bSuLC1JnyZrMmItxsk5Wc2cxekBrcvl3O5gXhIP/mQaNa9p
7fSkDiTAisYQ9uFAuamAxu/WcmJxqmqolyCdqRuI7tE835wJxMOPIk9ai4jcaE5Y
0zeK/dOBeHHvOMmWon6KDdAGY8b3OcMt9gxz9Hngph2ccbNXN6Q2Mnrto7E+hl9N
ThebRPDyXFBQ5qNmdJMBfoXVMzDkiXgzEQ4W6RA3UpMkJ4kZmxag9qGCbQeV/gGL
f6NCyGd71Tmk1pvd2ZYgOLjDUd2PoMj/K1qOPEsRd/5KUT3UMiK7L16viv05umai
JvwJ5NsFZJhYdtyk6kQgFaVjtRGbYLDh7fI3O36wxRJDtkP+I8wXladmmCFr8lHp
Hexz8iRNLHxN4FqoO33OTGwnt7nrmffpPsfrlW7gXGYAgyDzQhG9+jbvZxnIiDB0
NyDY2sSN3EIOvBT/8YrpvqQFd0g6t4oh/SgT5RoFl3ytvh4Xdw0txr0PmOP6tvJe
ZnqIGjaWtLKaEkFQUfG2bm7ldi4Y7T5+XLDoI3oWR1YIZvQcI7aPueWHe6d+T3D8
0KJNHy0RaQ1o02GgeMrVzyxe98PZLDQuhy3cMSy9yyTjv1kphGZKblnq4ejKnjbi
MdUUHyanFivx1yCCmEkXie7sxokxQBprua9c3xtQseVQRepIMMR2xroqkZGsuSUd
7cdCrfD7urRWFTQ1bZlALsCztyViLChXEa6jVNDUUed1QhNVM+cTQZRZLxBS222G
3NlQ2wkkBani58RL1EKrh1UbSr4VNmplDhrTKX8MgMjxoetZIpKC6bY+StaUK5kt
rjqR2RDahG5s+lFYfoSqa4QIMezLsj43gtSD8kNqY4gBfz1+oAIYItuYzaSvoDX+
F2uuvTVY/ZONMrRr0LTMuh8E0/C8JMePTeHlne7aUR3LUPMCM/lhtelF8ontv6G9
ccVqJevBm2NAmcK95JtLXSebf1DasAPLrg6urZxLiDHTiT/mhgnJC0TIVfqcQLGJ
IKrOKQDY2GZmtir69GIjtr/s65OKatKWScWtliYxXJgJBAinbYvgJpZAlvmH9vVS
9U8Mcn+NpJnt0TlJJag71DOGiOGsClgSHOtzFnFCTbsdOLnOcBUBpTjDqjbRuAbs
IV/gYhRQUuyh4qk9INLN6cUbUfZH61IYfriXM/f/nLyvOiDMQNvvEBavMbIZKkzg
HVqdX7zXxbX9Df1kFd8Jcl+HV1U61j/mfWE26vKfEYIt75Yeyt82oSLJrSkRubHL
NZf5lkBZzU5Lq2RT4v/LUlAEDv7IxoVu9dDPMmIZZ9bf43wumVNQ9/rkiYSSJ5dD
N/YKR9dCcpmZ9O/b0p6iomxiTcPJuVb2jaMl6tpntYXDHCpI2jWPmFButpuS7nR3
J0q/G2ab7x8S9gDZVAR/Hi4TfxlMeyp3nAnZh/vy6CN2EJUPt2n42KrySxIcIOyB
1v67UprNkGOX/J3XSwBWYO9q7pgRQEM6S2QK8p2G2zy9/OxnTruBKga+Ev2t4W6S
MlG456mPdlG99nyDCwoww4m4U3hB818fkynWOBFHyMA3WTU1lhkL5tJzspiWsRo9
mJNtM7S5B5guAYbNb2YSDTq6p1+NOKA84I3IrMvhXp4lIYjwB65kJSRMGF9Gb97M
qZVd3N+jUUE9dYwzGlaSoALbT9iAfx/BeIlVZeIpoaNu2BXhuELzbSHD5e0XAy9P
u+PGJzNW5w6dOEyjoo1vT7OzpzZATkOQryzWGktRseeBZtoHZMOb9wq61b7oTRan
1ZvnRqc2f5m45ySE80q6QpZFCeB5fykdHEmWWsAcrWmZNCAQeLmKajqBYATZ/LrK
doJMvQyTxUn++LfZc99lggyFyJxXq3AFvMSWL9CfqHeT1kqRTz/LHC2XPfiyGMW6
+bIQTWz7dveGQMUTmx4B6S7fds2hpemsXTjpPGlvc4BLEIRmbYw4FTW1pfDdPHxe
FPSIaOoHjyUSAP+g0/LHazgTl5+FebW3dw9pT1QDMFsIPhgs4+XV+xQhOcj2cyBK
O8g8PGuld8x/d+wFleBoYXWoSm0ptESwByRj0Sj963IYrT0dCkS3C+3cZIkhhFy1
cvYF7tSxsHbl60U/8IXpNKrZpV60qQAVLeisfZiwzVE8DwJcVG++FV0JXt5lydeP
1qSfW2m+zpVn+Cx64fWzJaT3RuDkA+uPHfYaU5B4rTFFShAwrmDJe1YC1ZJsJWBE
vadvX7JSAqXCmcdVmsxhoafrGX4KYvirL6oEkNMrYILbT41Nb/rOvxx2jFw/cqrh
iZzOs5CQDMg/w/jhrXwLMvpb/JXzsvyQZvmooerTYwE1J877872u6quNNNZsWeJs
pdKDy/zx6NluSgxBk6pQgLlz0/eR4cZTKx8rkPe/qPm5bLtdl2ad+Nt22bOrPBYs
2DKU/RnTBhqb28lclhewLwn/G5+7XK9F2zfgGrpPXX6Ux8cVusZXwiMHNaqMoxxf
rBnyr/p/ZM4bU3oych5oNIasuqMFKGOHb9pShcssNGnta1/dH65SB4IAciFMqIr9
dpe/8VgWcQcWxrtBMcVNKs4DKzPuurjgUvr63tMo+Dk0LY4Vey/ofdbikowx590w
1XLlAiSf5MI3L8BQ5Lc+38LZBQBMv6jnVQzr/R62sj7O8VcMKMiL8og7kabrHAix
P32I3VpgrpxcHdACwIWOvG7tOF2AoJCH1xlDzvnwwbSWoIWlEka3rn4l+ABpgO8h
oiKxrtrmTMtowHnMO+uB8aW1FGoYf80yZYrb1IvBXlZfJIWDIEMresKtV5qbMSAF
3Wr0tOfr7FwirwoO0MuIxxqc7hOUEgfNLD7g+pafhAaEEboBJx6cr8hgdk+RvN3j
pUwrMiXKhGrQiw7v/V59QvAmFT9r9f22EDXCpi6xbVE2R1yP9Z5iw5VQ9jZO+vr0
/eCXcWxHdIj/+M56JVo/XgeiQEdHEW6LHGF+fvKjeLN1ux5wPFYJfv11QTqRMdjy
H7PMnU2K60LhlkRg9w1BGPB8K+Hl1rR4b7Ux61jTb2v3nxgNyMiM/M5FZHEWpH/K
CrTm/6gcGu+ZkoJpC1Z6yDVAX8aoxn3weVmcExMDazgUp0OKL8Au0I4DmGmbrut5
XFFcLSejp25YG0wJ5HKda/lrYVQN8TiCQJ30Sm6u0sQJEE97x5xLOLgrfzSRgC5l
fyidg0eBiuwEDY/kMhrHIeihpd+l0Mi2dbSz2AtPjZY68deaHvYBnR5JPsxnR4dV
HkwIBQhSH6skTxk0RaVbbqSdWlUMm7rTDr5FoQzuDqW3UMiHGyD0hoGEc3N4IuGd
AHNzJ3IP/FZMV+ZzfriZOM5vAQbjSjVhRoyARtQt6LOQOuHWi/1PWIRXlUMjGtz+
jlGcWumP2XkIRpT/N08GbNEnVqoFujoi7IvNb2EDPoY6EBdF0Pts1bT7/a47uCN8
Duch0xFI1I5mvXjthkNYcaGev8MQt2gB0vMOGI01YwWJVvbeqNLYyvFmDBT5jwhz
5RVU3FYmN3TnLp78V068OKbdtDkbFP3NnDFFW/gKea39vEWsRME0torsyUS+mnK1
uw5TOFqffYv2rQ8pfcCC5gwFvHWg7dMoOOCoVgDTbaogij8iiRQmMQvnXLvhbTv+
eJ+wkRMTGjPlcXQiAXERQELOYu6pS5DUfjgotycqJbpnPxqRNVkp4w+jLXgV5PHe
APTQSqDyUn+TWXL0TCXRLYFTffqo0vJvkLDc2sn5EoP5MXxLLkwD2Ivwee51oIsY
lXv3t3Z/us2Wg8k4PZEUMaLCVeNvpb1qyK0mrE+vCjhzJasfigf1x4Rqz2OM3hiX
ssKGoAvQxB8O+im7mfGo27bBHlvKNtw4DZLMN+jzYJ2IvbVUFuITN/Jnko6yVCFX
QbbQP1mTWsIH01mvEvqVhx2Pe2myBf2NnuohyRbQV2vd5zBMcS9600/r8baw3x7e
7kkOUdF5BFCZE9B5KUhH1vwmO4Dtrc/rxIj7xCicdjha8ZIlppiJv4havOO5yX7r
gVbkSYDQ9gMD3ZsQiXrRcXjL8jPJgCe0DcwcVRAvu0TbWLO3ftB34OHkgrKiuKEJ
bJg1xC0MtiITqDb/0VTLKgx5z/Ufsd4GwRRHRapvSdEdbxkMs0tr+4pSRfbi/Xt4
GUcGj/xhwkvZ14Wwr3MDgXZ8lcMAaMlsHm6LLacHiO1AKLSMKOI9QLS2krrJZJ4I
wkNdOssox/dZCiom2pIaXW7fu3JOZepVj1DWdUivB16rODFgECEdT3wq+oe/Mw8q
bR4Jhc2rN6fL/6LciZ/GZftXxH9C0WEUxRp1xzeiL8JEvvODjv3XaBqtlmADhUJi
g9iFS2ij+Zx8XC+ou2+K+qQsIpP1OPDrQEZVKWFsbAtFAvJQ2BXZhAcZb2GL3saX
CQWf+BPHlFwh5zLm4zj3z9tIfkwiwVRIIHnMI06FJcjNtKskwrNKQ3+NiqqLpdKI
CziiEY8JVJ8i1I2gLDOguap1WjJAKRnXotqITsqFSJlj6kMnGa3YyTEBG/BlhCCq
BHsbmYmu0P7LEj9Rvkb/gS13wMieOzncGas5GQOAq6Zh5c/GucbmvEyx3xF+7G8O
Mr+9g2AWX55mCiH1NGmqFQc9DRlRIIEVeJ+l6sbNl2+sg4DQkoYRZGi0Y3c1iJGl
2B25nboIaVYEjDs3qWu/1fi48YfSZsu/KSOXN+JU6RoWHAWh7zRb4q8bi7Lu7+fV
gh3xG2dUdKy0YNtFajsLfZcI5d5gdK2fOQoSkMP5QkwFuEzPUum7rtX42tBXzw/R
k0WFlzouEleYX6zmERdBQsoV95FeuXlRByMdWZ2IeQ1fw78bfyYCFsStt5UIlLa5
cZczY+8TPBGKM3/mRFl/wqzZCWP2scKR/RTpVbgTdAi2+6mFZVgBXBbYiwGFMi6P
vbDNQitnx1Nn91fT8X76Kb3h/m/rOsDa+rKBpkNJTeH6XpY9Qt1AxFA9SV7v8WqN
IwimBfNk+Gg6WDbkbQxxQYpvQwea/UWwobO+NF0widQYk98pJH1lDk8B4I+flvOm
Hg0OG2cn4e6BCyIwZp/czDnsuuleLfqxGRe0UhhmF5pu6BJpFSLq7Vnv2SRosgwV
N7Ph5A3ZiHNSSJPGg5vz4rg8Q5jcZYNeltdf9TzD8ycL/0DwgFKuzmDqy1kgBD4R
cZH/30eJ/n2octzGHwrpjyBHAgIuz2/ABdscLwHNzXWpkl9umDi2KY9CKLJV8wLl
B/0H+eK//6pFKWNzMH7b/kZt+0nyVM/pTHxP/o9Vy68zYanxqw0Hpq271yD4eVil
sdCu6nYV1Z3M0blIZvQIuEnPV4dS36Ui6AVeti7itj3v/GoeNxSZfUMpHS7u5UzT
2yHyLMSLv8NibanNXOEXPYl35lilXfJaxCzH7VlFyI+erW5PL0SP5n7E/uGzmICL
w2AAOJX6GkBkr9zjcgnV+IodE2jdW9rg9jL3QAsNumavzR/+xvZm20w5JZD2v3qn
qns+VMQBWARQvE/2FiPB72Hk7DuNhSGiFnnae8Bbblr1lECdlQx3WLA1zxc8s8to
nq//ukKDQks4lQa+EJcBmDhs5aVP5OIeX/HApa1pw6yy1jDcQCjKOXK2XMAGo2YI
KsMzontGgRe6ZgGZKRYp78QeBrErciEEAQP8sPv1D35Kh/OjXCsjk0zGVmUeYoyw
9Zxv0O1JCslw9WJEDQaN/swCHjg1PrUJHsY5qm1HmzcuWnzOhfMbItDZy8setm/r
zLWRGOzIEy2qRY4unwf7LKeTy2W/wlhzI+ES8kf8glqKHQo20UyyHD/lCewx0ma+
WU5Xl17cB/SrtdQLUYcaF+Q7MWekzWkT9lFp8j1bIz0LeD/SiR743ooOqopX8nCe
mRluqwIfZRgv+vKmUVDGUHwyCz2n15La0rw8yWy5lkbsjiVYwNWa+bNCMBHMlacw
gOdoSXMU0t/Rp7uK936trIVRz+fmbQYZf4rkSXaKklCBwU4TAXNQzP3WBCeSMANE
vwHM9HYMNwDEhsX3D6gr4oMLhyXJjG96irOKHa+UYBBeAAb0H4LRHG8jZLey9Au7
k++x/hRkDmTMAMhrV1hmT1kQ18x0WLNdEiFCMpkyTHbf7CN0W9A1U3yHEm08zBsw
tt2rLK6UxabSjvS1HZBRyhZmBHYHF0pSPGcZfGjU++qyeNoEUdviC/NnQ8fnmeyE
TwoXG9fWmwGuDRF5J26BZiPMivZDSwOGH0SLXcs0kAH3O+VjSkc1mvAVvSx3IGGD
ObfStK9t0yBvVyfIqeg7X8PO5WOV8ARCEfx0A9RtOZ7MRgLSBW9n05CK4lagAKAJ
XOLKtjmRTiL5mCVkCYH2x1xRtqzp5/s2uxHL0j3JhePCJr3ZnekhGB15Nzwiy2nB
GdUP22U+vhohCeG6hf9unWxgv8tgmSr1p6gQDsLMiOdG5BnUBQs2OfcieNdY/Vpq
EAVTaSiHtYfIDrdS0a438uNF1VHZwiHidQBdi4/uvrLWCnpi6Uno2tMyWwLVp2kp
OiYU7LOx1vNbHiyYm39qytYWlV073a5jMS3BLYvvkeNtnGyhEY4RC2BcwI57XX8w
lQdteU1cGWHykFduOyxWQzMIgwJRFhdvrWiagtItP1eYjqAf0irHz9ECikzhPwKW
8ejaCFw/LLL/my+G8td+PcngkRwEfLgxA6gZNSCnSbMunOX5XB/SJPiTpR1/S+4B
Bxl1LG/IYmw21y68DP6zD3391hOk0owBX/ggIv2k69uS2cICLjFAHF1vQy8EFHHH
tEhjmQy+gTBB5E4rNMbHmjm/JRxSKk1yIyf3CQzLJIvFk9Wa+9xZh75w64Q3Avfp
qWrDPEKhC0mfYai5OVNlLKSW50/c0sv50qUKgeXUefmoUyWR8T+I1Yo5FLhyZnzC
7YqPWrmQp00pMEDxKAufeg0tKwhw5KwqbTF0eghMA/stXQQPRfZIPn/QQ21XDAYc
4uYjnz1JtAz37E0PKjbIlV5/NUqarm2g4uzelh0GaWOktvT25ex4bmoMxRomh7ZT
b0qzOrCBtfjbgxc4dAOEj9i1s5007YTauH0JuFdOQap3qy6fx6TdBFQaBgrd74Ii
99mzU9P9xRirvM1RAOwkR/usLw9ezyi0fd4Xzct8b1PJMWIeKxE9/BqutINtr3FW
Wuzr7kTkdcCxC/77zR6US2aPNaOq/c1ebOJQ/mnXQIIs6lsrlTsvGvHlFQRlVOgt
FRsK9goreERrBi5iRTnO++Dkq5m+iEGhnaqdLA0y5wUcSBdYHSTuT2OvIG4sST/r
WndFVmCqYr5EYPFdpuSQXVe7pLbYiZoh2ECVC/VemHMYX5NHJX3PQHih0KfgpMma
4ehL+CViWUD8r4QFslfE6juzAzSZJp0MT58ysYi/JE+ch0YCTXuJpyCJQLtuZKVs
pfaGdPxuRgFxJLKdYI5hA1nwQDGH8oPq1ucgCxPIzbV9kqGlxZOa5+XDGbCj7itq
qs1I7kuTd5eSZ5cq7pbXZrIsejdnnxghxtWl7kI5XywECl+PA/rP23Ta7QhSUVrT
hY3Z6CGpbJH+uysAuFxjrQbsTTC1dKTydwJVEewAXkmBB+Vo48g8+wyLga3ewPoj
EFpUrdwPMtdzyXjxBlz8qF7hUtdB/qbwpp4kD2QGpYEUCVYM6V5F0FEAjYg1Sr4P
TpajNBiCM4nq8QJQ8lIaE7RW2glJXVcH4IV3YaA+Zf/4r9T9eXL/xxO2P32PZOYa
7VmQuleRsrQlqgNkNPFIJgKc+zfjFxVXOwgrsk2Jkm9GykcL3zctkaaLoJxgZFaA
Vy8Vom/PMt8oqE3dNrvFfVimvMggDOivgnrAHOB0NPQDGTqVpGn74s7LFrWDayO9
Wz/IsbtiM57JEelfsovnpLrRZBRNYSZTYmMV3W+pXm8DnXDmNfuu8cZyrGNyT70S
WUMYLarsvC4Lb8SP3v4OedBh5X4hWPt1Kr5+jKU9SwNH90XTGJ001MxStqjwlNa1
YiFAnYMFXAhsZS6vPkeco60uYgtIMQcl8ALNPpKgg07kT7i6loWBZ/zI3lwj45or
C50pOnbTeu68Pi9xK3FtsPho+XzVG2iT2YbFAIw30ygr/oZNU+WzYfpV4KR2BS73
ymk8RpAdrp8I6WU2wCupV61E35szj+YYQDeB5HJKf+yvkLnn2Cd4YduOgVyVlYzj
iOC1gmMfm+u+C5xNHKkCow0f8i61vN7lNlk9Yg7qenfQZ0E008SkvHStG0AO8qKq
AlDab1kcZN4zOyCvQmV+1VoHh3t/e/27/gYn9f7yFWRoNzhu2GjEdcL1WXYjz+zL
1zXLYePZlgN9GWZTBL0MbaRB+Bz94+ZXj/SHiVr9WYHIab5WiWOw0u54PNfX/QHA
RrG1k+bGfO5+E/PxEDXDPZMRP/oeyFh8tbo3AVH3HBALaB+RvMYzNYc0LwaGphQ4
t2M3Bn+zyuzxTIwhcFVlM9U42a8FIdtnWIuNqFzgaJOwLT9dEK4l3H261tVmv5tv
RUtoxbZhlc2JMizHJSVV16mJSNzlwUrgaMqGCE+K67jahyl9zDBoF14uYoN18xTc
5seL0cHG0ML1iozVcdJCxce8cEOegZ5DB9bwGDgeqFIuYpHs4MHnYDJ/MsGCLB4I
45UfQckhCWJF2JcoYvRQGYAadhITesXS0UWjm/we10qJg3nvwjFLH5UuK/UU93wa
tscTl0X33ouPNIJqBm9bYhhfV+UlSaovXaW22boMcwR3PiW9AKVU0gC6vGLbe2IM
dYSrTPSk9oMN5dc+ZTyQwFYlZAF8c7oTAoJBuf+N0JbzkoSQP18lCtoC6OA/ZYYC
GJw0DaU5Zz0Usgz8GpwNa3V7xeGNTyzWrjxYn2L7/nSQC3IGl02YkLKWf7a3R/2f
BQBGDYDIs598vEiXwAOFJTY6LMpQhLO/1J110KC3FNlRG+PlGqnpo2Plo5WWVkIu
fJi9BiJVIwRW8edD5FcalRq2V19u3xoNbt5WsTO1XavTpyBFXVt/0pu2pKtdV/vh
+TQABp96ez08BiwFVRyfKxEVyTKgWxPA5lj8ubpp40p2wAWD/243sBK2rEO4DQvb
WECZ7zAUaLJtSNLLvgYm1oXAf0NCrCNfNCfsScysKyaht5bWSCaWsrczDokXl9oH
wh8IWOkYDB7asNKS8kSFwOQSCZ88cdGdYqzeVbSLzCSsYwvdQv5i6iEZ0dKcqFt0
w5N9uHA8wspqEztJ0GcFH+fyNPL2j/jDa+fuNoIlZAElDAoM62eZkRUckQCwX8y+
Kt+745ZEWQ2jXI3r//RYEWuXqlz8Bv5Rd+S0yRav5DBLP764+ZMVQZeS6ZZyFvPH
qMVeD19QUC6jXQLXPlhlsgc9pmijOQ2Y1x6kb/tzWfXTLZtiCxAuOG/OaP7Em3zI
77TcAmoy+Qzt/wwYM4s82Zg7BrK/8t+5GlkrGut0lmrWDBo1DBW7ZlZeCMRg8kg3
5+AKo9BqaQkePcOicSjPMffX71i9qtdAgwUiQUSQ8BdRTdzn9fu41dshFTD8I7B2
r/PkWvWijlc5XHZnqQGToxKTuSBsuFr2gW9ZVKr9uRlAgjW/6J69JtR3o6zvi2Fr
Ds00nEWHcRtcAV4o0B4tMdXijiOk8oBFjTxqqyCzREIMkMKcX8GXEQPAuH7cH05P
Dvl1IoeEXG6KMZrJ0XJ/7sXiLHWwWFqvSSDUO0chCzap7/C0HK6UC/qeRGI/FGlR
Ei9xNrgmwUrxOuLqUhNRoO8gZ8oHOQ1oZ7wBuYwWotvln4t92pG3x/w5/kct3SuZ
zofXiU35NJteeuRyxzCxPMz98BO7ays8IdGsvaghY1rmdmpU8qnXd+Fb/dWEhFJ1
6UWK7T9BDDh3FEukOFQdHPFgQTC1RcwgcHOePjWDyLBshOvWKUqwQ6UxkBMcCOxI
oRFfoK76LWti+pWLm/Vwr+V/fzFc3O+pNRxBAeja2tJ63LCwWR2ZkQgtXoKhClR7
Oh31qrUE0eoNULV7iQ7BFOyQsWw7pbI7E4sbDPU94UZH88MrbLUEEGAAbTfHBnuw
7/Hp8eE8gXuO4dQbeTHlEm2s9kuvHVWf6C2sbNzAmf6q+IjXN75XPNtgWuDGeaUC
P7WCORp07VgeC6tdv2AQJUgoHa4yUTzb7fQcDOoYZpW5kLXI5OIZf7ypRNo0GgHA
IMoH5ncnlzZ2fOcSh4gIpt5OKYdl6V7tl5XOHFmqj0Di6R4YUiKbsBsVeDNyq2Aa
lekNrkeB2RqCnx+epy1vNq5ftNrTUVkKIp/sJzP7wJL3R1qu3AZ6DXFf5qxFmEmQ
neWRETsIEe3SShnbrby92sgmxuYNWZZzBi06a+vvuC4e5Uf9s5GJn5l8nTdp8V8t
lBPmBxbZvO7dLiNiiiGCs1If5GfPF6MdfhyAflCR6Me4jxoE3bIy5NhbeJ+ptfBm
dcG5sO49JSnF9rbTEHe0HVXFdHtCvbqLVm7CmGkmeJjUzmbI4Iy0oaF7eU0r9yho
BLpthHW6iOV42CycyjxxxwZ17WuNnk/twBpdrvCXDU7kaUw9S/zdWn0n/L4hCVKG
s89ZwCIX6phT8PKmcA386XWOCEza0pqildHlN9rnM4lCuOIgHmsjU2E7eDCjUEIL
6ECZ+OaqLyqW7F1GRY1b/B+ZJAGz/gugZrnsqqvqSxI2385+EqHJo80SM9OfsPkt
D62kDkVyqI7h+DxOkq1LY4lmuU+SsFi0mayyCPJi4SaRkBwznQcqekNg6FX2cF0b
ukw0g5M+1xXzLFmP0UkdrwFecVHUw9Be42VW8KBEDcDbRMHJxj42S75DZfxJu2RN
YzOS+BzhcUIwls3MNEqtO+buCjNquq4fff6n1u5TULwOF7xt9akeu4ThJxNo+fam
LubBdJedxc6qBWIpWOzU79G7PSY9Kx8wJxg1qQv7eU3hGZnNSLFEY6GOwxMiqM42
pW7vSEcrMclCfu/ViM7jVwLLlKbyTXl9T3dxoNYDG/+0FRhBepDZ/w++J+T8N0E8
CkssjBJD3BrMkGO5okeIXmKRLTMZ99VYgqK1Ap05gCXoxaiBDZv7RQ9F3w0789hK
FFh3NdXLiapCE7QiC05XBas8hsPndbXdtjQtnW0irZw+r2pjbtHZVpya3SzyUaTI
nAysjtpCu1iTAZkuR+R9mTVvCUQ/a5+T8oQ30lWLYxOdkdTHo5LWK28MNUki/7Vy
Tp3Rs5r9GrWNq1QNMMCXFCGIxzq2RyyJH2Y8s7p9TPI07gAH76UBArriYySL8byP
tA1ei5XIIbUUXpu8sdtTG2oqoRUB3Z5s9Nh0z9VMX+in7iid/a1SobH+yvm2n2Yw
NEbA4zaAR12/SoOent+EY8NiSYNk5J9zyr58olxxHXthzjlK9NctyRtFAhg0RXef
low+pMeDrApapOMLbb+giyz29vjhkSICMasjSr+lvwEA06GcLB53BdAqo5M7+EjV
gQ3AHkxunp/h7ZXnDlm5xNYBbV03cfAnihZGiVZFdnvKVOEV6VJZ6UvwxW4zrGDn
ckBoTu134tyeOIRfpzHBiBUTJCVTDal4vngSZve9nB0UagTI2I4wNKaTLseqP2j+
co/2m49GsVdjQN7btYtLdAdeGuhoAqNmKfQi5IWWqqDm5Loc6E/Z6x5iUHUGa3dB
iBjmDK34A6WPvNzzR3T8C03GrQt4y31YCymcdF1K7Q89G28VyNEaV/hNYYCAvYmL
MvRGDbBXokSbgh68xm7wBcN2DqIenKKb1QBCWv2R/E1PlGxD6bazfbJvmlEeyXJm
UaA6Fca8L/ITjzC+1UaUaCA4L29PKNNHP46gfL9ivBX7d5YSD6KV0BV/5KrDBlze
S+z+ldOuXJSyDeIGUi/TjHlR5unGelIBa2n7MblbNu9oECSY3OF0vGuCTW8saKSq
xbfS1VN+CxgWAqYlCn43wEXSa0kksJEwPgg960/zxmP7J7CU8dkyBFCoVW+1PPbC
m8IBGvneEzPm8sdQYsWFSUuCQp01EJMyZ/npjAsMkB/henn/cEHgnLF3DIak3x6l
xrKbbd+/GhNWAW5lhAJiyWrKnWbG3KEqkP8v6sj0y+lLssbh6V7iNmbE8K7GvDh3
xyzIpqfyL4FjrskSwnslYuC0HWw7nOCL077161QZfaVMR8GJhJn7kOb4inMGhw/v
TfkvYo0U0h2VqqH7enH8hldO5C7T/T6q2qBnTr2rsjWuU8wu21ecfIjI17NLL8Zr
VH5CU5c6I5CsWGviWuK2A5YR1/TyEwQDw1w7VU92812n2Mhg7EbdLS0QWfj3o6Jt
lnzXHXM9jnj+258sNkvsqW1L7yXYlyejohc1UHw/w/XUB2wIXEG8Cu5LEAyy8EgB
DOGa8UQbZeQmBymh2O3pUIG3K1VZNWTY0my77jRLly4u1juyp/IkSO87IoRyCE3T
F2iqYlqwbOIkkscufwi/LupKWOlvXTc+oU1zfC3nArXwztvnwznfldEEIFaWw6XP
OjENbpfxqHdTCYPdqEdIwSt/TlaevJEGmFZgspaICzjmdB0Yws2KdZjeMX+1is1U
q4aAxq/xo6jQz/rQRBBiE01IOHU/mgKsdqO8tt3lsI/uorhb7gOW5si/ktwfNB8a
FHDqPpUzKuRrCkty06+G2zIHQl4Hp30EUwD6twbzWZZsjQ5SiykQqvbuQQKh4j/8
pVIdVLadr5nUmeJ1JgeoBF4N/MZT6ulji9at7LNKqHJY5g4ermPleWqDoBAFdQFH
gS74lrUFIamj3woGNIX8hj8h927Hnqx7+A6U4Elz/hZCy/MmtY/rXYcqeeWpKgml
KREZMepXcIoBW1FU+nJCKN9fGz4FRlWj8gZWir/QzcEzJyQuCshX1bcrw0mNCGoK
hOZBhd9Rm+KNsz+OPY5bHHVxCTePes2ZWfKaBoCeo7R63v0BZWfil6ooZ27o1F5w
O0kInpLe7AcbekYP7m13S/YRur442oPOE4TZ0UPpyLA0g1TniwFXeU/C6Zr3fwj9
8V5+hiRgh71Pkx7J3vkTZoyycRDwoCkUUFgJdrBAd8l8wQYO4z+e+VYrxAoS4OGS
7EOhjulKC7rUJgr0wTvkmcL5kRs5T6oysJ5DhqcBTFBWmv/ySG7agJW846eULmMp
hqiCpXnU4Id50lGxqhRAKkxULGB3rk9ARBlar2Rr+hL7PItCZTHG8fNOxBZy7dyI
SL444yL9yHCKhT5b7u0JvoHwZmLB9fvhwXa/OkNFmj0yzq8DneNBmZPr6d51XPE4
9vw5TL80lESSelgKL5TB4FVLdGHcj2HeckiuDPB5N+w19/A86Gc+H6Cc6CVw8WNH
dA6A7ghzoUyZrvT8ms0n3jZrXDLL939HfhB2phWKbfP/Z7AoqBE1iSd7KDwL+CWg
ALdVKUuEtoaKGho+kvDplEyGJsm3QAIrdv637WkBjmLY3Ifpwpjfwh3cgz1W7A++
H7xsXHUZgfVh2TGM8mb8fReP9ftKYNQCos65OmEspuVy0JOX/p8pnm72oBPI8NMF
IKzaGsXmeaXqU71bFeGRHTgSVBGD/uMbNKwX2u76tDNUiomN8LspNF6rs6eQ0Wlj
+PBs32cQtywU4NRYLNgVlGFY5L+MOox+v/w8kT4YjPNEO2EkwM0OL0Rs697Rggl8
GxHmNZU1CBtg30iAfo8rT76WD6172Oh74/Sgd+8biCEm9si1+X1//qY8eLQ0mVTr
aqjAOmlnTffcvSwK24MIbvjHO8VkFnCEqx4XW95DVlakQ88yVsiS1udIjjHm8YOz
I45uiiXQq9xY93qGO8Ajrpqsi5LwWzYoseVqPIJLiyGJK/01ekPHyWSdgov4kXJm
+NhJhNAK1GdDi4PkeLGOiifu8V7sHxpBjK1N3nahEcQIdDAUrXfjG0aDbBj54Typ
CqqRYLBhztw00IssVW6lj6qHvGU3BYhStVynj5TTWWCrLNH0SW5ttaRX8HYexVRL
BX6zzpfhJSLWzEMMZfqBSJaZuE4m4UBzRxBQpnu7M9IZj2gej5zLfjTeQMuRXQEn
ReSMJtP+xGids1Ww22fN0icdTsBKfBtlTmaTILV06duf4KzXrOkjp8c2E+yltLF0
Mh3/CWSOdgvZlUq10FrBplPckfNuC23rSnvPvytdj3OOTJ4muoO+KdSeV2YXr5N2
qR+c8+05MRu0vHOhc7p80bhT/+DBpA4a28/VV+mI2WFUUDPMm6sfV9MLt8GsyfmK
ulCCur6KSujVbSPYvEKrIxpGKgEbzVytSEXBuixkkCxqL9pth+1LMWYV8WvpMsjo
2GWegqhVoISFYio7IYhXAB3NB9F5Fa+51HXQZGqpaY33qJtohf53FsNjqBC183SY
HrHN54VSrEuksAPAQPR99Sf26yWInXOVM0EK2eURGHGMQUcIKRygrM1lVS6wUdfX
XD9Id9D2YYd/12AaORwn3fs6oVfcmL2z+iXJ4u547g7ulj/YsvRgfIkUm0tVuiUV
OisaOUZm3U1cDS5CAyzKdSN9agUD9DBva/0x90Gz2B5166Wfq8xnVwr0IAPUEdGw
FlXjPX4znwDaFa+ihvb9PyyB9gG3K9ZiyKQfUVw5IcIDEn7SjJbweF2Dzd1TbetY
CeQxy6tPUS/MXyJTObKlpnVw9/6rBVm/rlNZrPS6KPmID1J7fvuMFMPerKhh0c/T
3+CD3iGx8ILQ7byxmB2j8P+DDPcVUxYo3Ocj6Kb/pD0JF9TxklPcQ4p1KQyc+k+S
yc+8IuxGv5rnCRow9dz2h3YBmjdc3NCN+Y/FSpbqzv5yDHnh/4ocBdAMLoymp9i7
O8YXxuwEIe8QpqO7IUmTnPD83JeDJJyUlTcfZnazRWQL39j4pWwUvRyc7XIMeXqD
oHs+nPkieM3aJ55CV4nebfiJye71RKe38PbPX7D8q+3h1t/+qsqaQbMg9QMK3d2z
nTLjqlus5C9BtmDZ0VK5Veb8E/GKNYkiSCoa6fZl8vTFlLCAiDiazYYpgn0ykrDB
v4wfdNHST8sBP+GUmWP3cfl7DBkE0+FyxYE9wJfXu290GUPNBRRWtS37t5DTpDdf
DKf2f+es7o5o/8mqXb+4mlLouG72+jRHyL1uA551CvEbExPglFMK5otWphBJQQz0
kYjYi8NpZSUinWWHfqP4Q6eovZOPapUalf8xcVq0tBhh37ssK4TtlsrwO1G1BiRl
yqSe41+dz8ZcSipR9mk9MlGjRrgYMjFYu/A3yxCmmtwnr1x+opRht5XF09EpZgPj
cLtIFfKdw85OajOqXW8tLgVAt8pEDkbTCmYXYU0Z+u0y6/vMBTZb/lPEq4bs1EPp
cREefV3pQSKefX9nOBfbZrYUt/vglMXkXz/JjwO2zofUaUSJ+A1f7PSn05tsRFhJ
rjQLGp81AZ7QPl9bJb2T+MI/p2V4OuQmQ1iEOEdceFSSq7QV5333hDqb/DD6apCV
WWuY/1bkOf+gECgOadSAEbcJ3htovUfq7X6WiD9L78qGzajjIqXCc04xuqlEHP+3
q3mTMkEzwbheIgpAQhWUXw4RvX9uhySccJOQN8ekwH/xm1ZAwIwp0P8I11JzQBYi
v2PfFt8QIB9JuU+5cMIPCxGMu8ZSQGZ1kxxATZUMT+bnQ9Cxf4X6n6SwprGsY/hU
gt5lfngrCcVKtpYqgZgZps/oChD09KIK4gxWAxz6spXpX0sFIdbBexK2T6cXlWLm
Y9gP85HmTvvGoS714jpIMWEORl7HzUQSGXMoemCoGMgvb8E71GNWA8wrZR1/5wcq
MYnwcsvDd6pf7LdWlo7goeD2JzCn8GHB9TViW+6ZY4ETUoxpXbCmjWadwbWH++HG
C9KmPe2uo43P/To6ZL5OUWeeJJxCJ3FZIdT0sImbF5/e2NtRfoXMRy3SoGEdSibk
nil0qG5uXz29sjmBFKN/FyDXx+0s62r9xGZj4zcPa7BW2/pyXft8Qp+SVN+kEgyx
jW+AstXGhlDTdswrnu723hqIN80SNQVjWoXClksZektWV2APepRWR9sNn0E/vGhl
HJbMiVnJMqP26wedmdyJqa6g04IA6XbCSqh0felSUQztvI3jmLTP2yfqObnE08pO
hxt4RiHK/lOIzdgotSZjlL0YMVzq1AJJUzz2TEUgH7ZfZvI4D/obBMZIGr9cFj1e
87PqZQZdamKyPfmSJkZIn+U1yAdS1JW1ldcwKOnkZfgAiOp+rZek3uoUkfZSXiHT
eC5pQc4W1CNQ9o4iFNBI95wAvhOmOhIQ/dktotRyIsL5qu0qK0s6TlKtAkXNvoKv
5CItEpsiRN1chRmsnvAPHOFkVGS9YU2sgx4jR9QfdIQa6paxc5rz8SU/9EoHKhEd
gx6m8krD6yRfrHzPlhtCBeFVqvrKI97mhHB2PuNJWDyiJrvLP1EGPRKKcs69oVz+
2sMt9PCzoAkljuRHVLK6X03nuo7jmSUIcYslklbg3NPseAkNSpaBmFRv9WPLNFyM
vxDeFbbEebORLHWAYbDXOrlNPl63xNzhw76tqE3hcslFe71zrNwBGSF9WgPmcYfq
5IbMDOqXHNOsptyrYhZZiW/BtKwqMhhy4c0XYBs+Q/yDi2Bk6pYlTVDoVKOH2/MV
aOhE4rlCTFLyxxgtlwq4M2YLhFPFvcOp3oh1l1xsEVnOAQeiPOKms7S6oExx8I9X
ErDmUTH6JgnXkuAMUwSlS0X7quaBZuFpD969Es3vL5N6aw6iFuDl+GAFn07GgpzL
6OorVj5cbrO2pWnKOF2TJRu1qp/JnjWV7hLR2sUNo5SCTnPrgenezus09UVLaq5m
nm8fnTNK4ch3EML1zGIRSV1OtinihdzJxX+IOHyqw8cdKXv2t0BFBWv1LYXlW+Gu
FfszsrpsLo/3ymOWUsU78arR3aHQVSekjHR/GqZrJ+U1XZkElGpt+gQJyqW8xBS+
UsruBqdniPzfItLmKVv1vF1Zp6JFaiOlUjnW0TbU1wWPjiya5DPmafDX1C832nYq
HLMhQOgoonGT9kqTNICW8WqIpj4NX08DhwBUTEb90UjawchIH7sv/7i5tpBj7q0i
QWlvI6q9YR1iwhH8X6QP2ToRZZZyXlwI1/kF2zwiTK1GHP9chyXqu1dzbKaZyf4Y
hYOlhvIAPlEmjtra9V7QsDHOywsY6++yEtUCylB10Ke/sFT9LhPsC5rH4Avocuff
tzkDqfhvG/pGPlM0/EwiTP6sfQ1MhL/ObZgdVJaCeQvUcAuKL+KKvJW1EB2Yycba
23g75/+zsbF9AJlY6UhuwwF2/V/IXp+sUObZA9rGOaV8h1XKPoQdBbanIP61PPms
2sHWJh5EGAmBnxgx5dQJiB+xtcugqppUaJ3z7BXpV9vbpknZzblj2XFqwtUeHQLB
vnX9rfm4g90rWqEwzLr19p849EduSQijvCdwBCgTaPQACPrkh5TIFEh7wLT2jdLg
a+N0Mo61TqJUjigUD6jhCk67p38qyoAPe2CrWmhGfxBN1WLz98RKMLadii7wPr+0
1yqYQJ5Gi5YZRba4UO3MiBk345scww6W3yY7A4sN3G1V4uNPLu5WzZC1X+5Ya90H
vH3W34y+UbrpsJU9N4Mf4+avG6NKr/TouAbgtNZmWEf5You3MtXfILXcKx8aOOVu
f+m8D9BtmNui1NY7K065HLMf930zZqkCV9pK7RLjHCil4chhNXShtUz9IX6qEj9C
gnZLvR6qQseGQfe3G6mAjiCOjrAq4kWFb+wrsqltxqtvGfxsKZdSl5KVAk47J4zq
8ndNUaBpX7MN1AhX7u9GlVHF0Ls87BA1o6wgWRjLVukwX3VDJEqgurBMhHiOyUkS
kc8F4gc1AU2mfv04RLDTvO2szl0WUj9/Ho/Hsav2wPPsN52Nq1D08VgYTvVOq/he
hLEdQHqVvPzDVboK2GYLyYBQSgJmHgQLw7JkxircdG+33X1UcnbRV5gwzMFfdiop
MxnAnbG2QTjtkuCTAHbVu93mR6/T31qtnSDjhS7pjPGlaNLsEUmK96gxuF1YuqLs
zIcsTmE9onq+KLAh7cM70U/Z6u+zXobxiNN+E7nQdUu/mMddrFEqJM+YY5CPQZ5G
BrLS5KeiYHSL88QraA2ekKv+MneKWGhNM9oX7AOToyJoP3GuK1eyQrIxDIO/xw8l
VtAT3tTl86tBBRlRQbmFWp4N2ICGKeXQSC84BudeUUuGQt2sJaes7X2xkp0kpL9d
FIwuf1m+oOnCG8U8aFg9J2HmXqLbWBVycgql0SgTpr1Ue9othuFjqKPLpGQfKuAa
W4Eis7Zn8tHcAAMIhN21RtLt9SwGqe47iNI9FK5BF3vSPnPszLrpNaAXomxjb/xI
1mgVkv4IDLbYrU9Wcq8KmjoihykdjzvU8v5dvyb6ebPQD+nfhkXlTPYnqP+sUNYc
H57YV/FNN2p4o/n/RhlSPu2Qg2NZXbCzrvCiP/CxBoJaukNHdQV80YjsVO4nbIan
kOg1LPDUdN6d1FrrRCm4unLVDpIJb0scHU2n8DeMvBUYjMWQA1euXfxgez40TAb6
Qs7auAEPmO6w9noZLab5QJGt66RJmDPIyiJRysNnbJjAdHW6NDIFo4S0mSqsQtXd
o2QiqaT0dHCiHXQzB2No4wXlQUmjv5y1vhF83DMuYqOuljG2qDtnwPUk4SVXHZx7
DNY4VA3CPLum8iEJuiLPaEsF6Y8XgEb0WfQcIDAfP/sfGTt02TzRAMu0BNl5q0O1
sBGHu+ne1B49Q/3pHK9OZOckFxhvlHGpMKaJxTZv+oLxuyVdEBqlniPKpgtmPh3I
MEJGg6w8x5NpMmrWOkvJ376UAQGj/UW2EUKgg9V8YaNhIbw8QUSP1nrqNl5fjkMV
rn8ecTpdjIqjOHdJZ1i4YfbynIszT35ETRAGIbPWu6Pz84gjAFkHdXjkgCH0r0oA
YhDN7k1mVXH6C5/6lw90fvjgAcVzJd+NHSfZw/YxxHqTBhd2gd14tdv8FNHS9lpy
sgK/fnAGHwwyBqqocT0R9aSZyxq+DBGESY7sJN6B155hAihLWy8SrUvWOWb49AtR
diWK4o9srITY74jBItV5eOdaj10mkSUptA10P+LI7k20B5/MtfQVZcPCFa+QioBR
tI+wz1tMaWkiwr2masn0DxtqA+qp7sGiKV8vjB4bZ3SOCX2t0rbPA+BvQUfdUq2Z
zOnSB7Liqvz1PGzKMPi5Xcr8y+EnPVshMVmy0gYbWifB94py3q3vXY/m8WIIW/iC
gFcfa+k6H97kXHixCsM436qkN1BUD+dCZg3IAAGq0ovYOVc6nsJon387ePWQrgsq
EoqEyZW9PwuvjMMkALy4cYBAiGBkTwYlE+c5+c3u4TQYtQsms1tr9Lc5kfE9+2bm
YNcGrJmWAgEH3PyyGWdDXcVYii+NxYxwm0f2boBjgpwt6uAXUHZrBTCCWdDbY9Xm
gt/OBIb97dPT0CFFPZMOzlUK64bZ/T05Q2C/BMzq/xO5LIibYvM/JhDPzJYyHN/E
Vu0ucYLtbWXw5Zb45hosfoBwwb5yMV9MoD7KKNde2rY5slEjQPIiXH0vJV89T13G
bF/Wh8rfhXsbaZRpNtuaAanMx4ggUFffJlLmPch/ZlCPwMEMp4Ci50UN7f3fYF8N
xdig3paxhNaZpBm0AT+Yjcl10JuYW8BJecGzbnNIp32u4/rmWxbLcuY4GLzn3KXO
nPNRx07GYkjishRpM8u4KTYcqP67szRrLiGur65SW1i9MLRX380Dhx9ubyD2wrjv
gk+SPjqOXFLPmYtORfP1E7C9/wrnakIdcEmvPVhPq68vC3spjXqaLKJO6E+9CtaB
Ne3dsD8bW2hZmHBx0qPWIfJRMKiaAj7KX4t5AsTvbGgjw/fFjOhcDfmHdefskcel
/voIAky/okJkZ9LflWVtnVkI7GMaKR7JMWlVb6YmmheOKqMnkuVhgfgeTH7cy0U0
KxTOg8iFGUQgtxeQZQ/4kidJnZhowI67jGJNfoZwNrw5Sj0Bqdi+8pQAK/iT99UP
I6TTRfJTnvfQCdssFFyr3xomnfYizejHwYSL0rDARngFPavDmR+cjy6Ljnx/es0q
Gw742BHuGRezlFGXiJiXWnsTpB+XERkoKoPVLUD4ctXFCTMv3dMIN7w+yndoAIsm
XJBfe5isj+tR38xeNG2MJwsJ4dkq/Sh5pSW2Um/yTA1cQ1Gcj4vT9Pj2aJV7n7Ex
+/A1Yuj2RULVHUef3f3IpkiWkVoUNsaqKiL7y6Ajv/aWZP9W+rMUSTa75isPCNHq
xPfrbZs1FlGsP/KUu/sXMRCx5KiotmtCHyLWZu1VQgjCmLvAz3rEnYF+80cq5QqN
CRySAAgO+/zYQGuvWBQzoJZZc9BwYvAu8QP+DW6K8JTuD76zWG3oMvTlDDLN9x6x
JUPI1oKJRJ9WeTIyj/qZafGZF/gYccxkwK1nHnaPBRNFJrmAlbv6mBHDXZ2EXM/c
9bI3iwdQSL02tha5OTbPBX4QDMX9bK4Lu6kAI7Db7kvkdInh2tWrZwzL1UA74eF+
Wh2z79GmTBj1Ayar2dctUDnKsl2wJMNmikwenuJ2iean+qDpDlvlEssMqB8nOOjS
I8WzfmP32WHqChKsz9E17vk+ae/UDLODBMaiZkqmG/MCoujErc6UBydhBRCtr+nX
YQKCbb84rKSWszWbMcf2WFZpEE2t3CZ0JWjboFIIUBBw9l5EKwyIy2ducWyvLb6R
yjeJwr0yXhO5RYvskFqjfSOslUD6fEx6XsalmQbeFNkgblpF7S7f7kRG95TEuy09
uNdercp6CYimmzJD7G88v4rHWgjzVhQmx+9Kvd8sQOanDZdGfPmHmHLg8gxh0qgm
FWeyq0j1fSoW4ZUBA32a9+pRgEAr4Xm5Uf+Jih1pqNFj1mGIvNgdMvIAhmMo5Qgk
IsaGU98XbVewZtvJAbzdthBHnO88lOL4Anu7/N2N7l5dFPTk6Hwg6vdSDnDsHHBg
czpIKiFLQg09m0EgXvuDyfaXvG1DDY7/D126WODrFOy5/sPuqNvMLUC6pJvbyo4w
jwIS5OkcFthwiSQIlggsGUbmMHQcUsfG8GjukDlw1HkUAgBXec4mi30Vi/u5luXx
0y+EjeDqiSq/Ik6qruVqenGr4otySf/jr1rnMR6Ae3sP4otZCI9sTka3le1QDplg
+WMyZc9HGkyCrUJw+LQMb2x4g+bCmWIfS608FeUTkzYe9bewvGeOzJGHQjfWXRqX
8N4F1pz7HV0Jw705w4HA0e1EmDDFG74MZJ/dSkTd18Wgf0xfjlk3n9jJRgzwTgSL
xyKZbUOABHz7h4xdMvAqTzUztiCFYo48Em2wo1L8PgtG55rWdaqVODa3wH3DeN0L
Uwi53looAQGsR3vyYqWn5SFfavwfcYlQ0H/juv6nSt9xtKFsPz4MtIY1hYjZdvGB
fC96wPAiWU3n0r/2dTnz686bfrtpX35nLlq7DgHCcCHEUE1+NRwNBXrSQlmmuerI
CbV1kKABQeIueQKbl7xngplTYjmiC7PAfSifCYHaWV3RCYnBgthAssk6Hs0aDS+P
52PeEPvNBWyHOdXs+tXizRU0WBrRvywi8wqQrqYlwhpYMCrGHw/d/5wvls3vKLqg
lT/H84kuDEfqe2u7KTGqH7lIMkO7Jyrwvq7HmrqL3TtfqW10c/Q4Gh5GeVcCN6Tu
EHB23GVzfSNapEInXfcppSU4aHc4Tb0zgD+RlR2+b5TBYKX5ek9unHIDct/Cak5Z
8qmbLqtD/lOF7m9ipNodo0ExrhKJZNzGLY462oZBpEU6Enmp5lkB5oi6LcL7eRXK
yVsnlNAIAcDoB+wZxcGM0C3J4IuuT5/F7IS/1uLkZpPrb7tDFmiB/e9czRrHTWoH
420EucfcVPIhFirmeTqqsVHQeSUgNIqjFqab7K1W56Rj01phYbhexfOJpMfeSq/B
MPb5cXDJxLh3G4CvOFMimngQIR3z5v3Gn3UGHSFzrivtTDByBSF77wHvLJsV8/pf
m18Y10jXJtlK6DAut8K/15Qa5eYlQTY7FTa5qE9CaRXB1UaHUbg3xyOI45gu8CSu
foMz2qcPtdVktga23CcP1QbyM+qgdqVpJ43laAVZmhqkQ3kr5o0Ui7oR5/q283uW
XHEntMc1ZrPMmqSyYfSFIgA72ixfkH9hi5STf23ceP3m/c+daKjXK3FMxhOR+QBo
1eFFtJ8ZQ3OfYzpuqrW4AefuI09JOWxHjBs5rU3M6kO5G7SQ3uw+82+V/gfK+xtA
i1JUIn2lXybfZjs24D2mpITFi6VIKyZ27WV/QCxPcFwKvc6tzz8ASt5MfARCIiei
R34k5b862C1piqUrQfLWrQ601IPCeKKtKa/ZZoxSOyFLJYGBZHB7z2Em+mf70/44
U5fdgPshU6roxA7wggGi6nRTjthbSCW+FUlAFdYz74hvS30P3hts5AO9MmEchQqe
v1AS+w2rwALxWmkIQdTguB39lj3ZjBYXpGF+BYXaCAFQqMJbJinuCnphFGIcuRPq
LMfU7rrA5cT8DCZVoW4RQaD4VanRlI25LD2DF9rTZe1ABI3jcmRr4bB/kbHe/Qwn
yqNwzlETwWv2YRnMnGpN3+wVCbXOrAbC9NU2qQ227jHLjDlVDV0ENd+vb6nM0hW5
+tMA5dnFFrRw+wYklkjRoQW2Do0W8fdvCjeJjfZNJO6HeweAj9GN6dT/a7O7KVBW
aJaAereZRtJedjWkKVGU/FQWm7tjxjxKVYD4Qpu3nnq3t/CNZ+oHoI07yHjxKx7F
H5xNPYPZp+amcyc8agIZu2ftSjZDyP5avHgkjIWuFLABlaR3QbRPE9K9jIj/uDbi
xs8Vxd19mm/lnbIH2SlLviLG+pPmG0740XSk9ZPMFRqIL2V9wrFBbEKjMfF9XZNM
kxXJxOewnOFdQz1/TtdOH8qU8xUo8p0Dv64wL+kMRTG5yaTM8xoZFBxIO27vX0Q0
6ropqhbFOOXgMjTwCbVwJsYOJOpp+OPOcr7T2FGQTELeGLfPoJv1mUiYDF+Mwshf
dMR3SPoryZ3Fe9DcTT6AbeG4wtyglLMHfVxKP1wH4S3DGz/ni++yMNIsWzmUdY5E
Uh0libhMcl2bQDbK7hgcCHUAAVnn/dK8czDmSxv/mRRBgsYBMgMzHao9sGqyWIEP
6EGIPepaqdiHD4elSYCV+ZqhhDk1SPWdpxgnqTZA86+VIbpGo4UAl4wqNGbC7Xf2
vBX4PqCg3TWyv4SoXNSrz7t75NEDSBpSbMSs2CuHdClaSjSQIrkcrtlcoC8HTfY+
evMzfwtswOLTkfHYkqbr5rgco8AYowJEKkBM5dlNw4NjBasc8Ofl1ScGKguwI+A4
Kq2c4jiorYeIflonSKsEHknhchAXBMhX4nFz/jZl9pymO6tcrzDnUUkPQdXNyOe1
O3Du2jAyYNGjeop4fsJQNsWQ52O3exyG9Ewhu8XknmjXpt4CLgH/YBYGQAQbT/yy
fmHz9lQ3Ev7yWjLwnAPzgJ8WKnKg2JumRG5oCxYeAJcyPk1HZWeFnlSUTPxtmnqP
c2vq6wvBFUdIyX48VVL0eZQmWWKCCVSLUzkZNqBoteFWuvmdvkqtrA+9ZD4riR86
4Bwl+oI2adszva1dGTRJyT1sbMjo4aDZxpYw1E5SueeWqQVbN/9VcR1p85SPwbwU
l8bQN4aJTF7V9hID5IIXqRwQidALliBIVIVlPqXu687Bh7+IvJ6F8ihgiEn9j+aM
ksDzd2lezOlmyMsqESn6HQrHGrpjHDijKCCWU7HdJiX7WVcg5Dz2E7xM63kIsXo2
L6sM9NQOiCHox2YkZ6HoBqlipvcLAfwnUGAxBhH1CTm80c5x1An06j045PM0gcXQ
/x0mI7Se3AD3nd8XFsaMnSlfXjR5vGgsEqNdBDJc9Em3OolKMORjCx933gvLMbCf
zXp8n0FLjK2oqs62MdZYA2XnSIGExINk5uOC7lJ2wh8fXwJL9AVUtCp2rdmn+/Xm
TyJNahmKnCLR0KaOJ2tw9EIDoesejgx6grCN+A2G6At0gyy+aVx48horI2af7hg1
YgbyCX3MIuYBgB+6AfmJN6pKaj7VLvihe1VNsTtmVYLj7KeshuSCmC59d+Zrspq7
aJQv7xTRuUx4aTvepfdW9Oid3GYjU34C0YBc+4AbWHyaSpFUaArAAXx8ddaZdlWw
db653mpdBvTOMRAc93JVk9htc20PiC7++6X0Ys194zhAhdSHXospDF/aHbMitVm+
4bTjzJMegBLjud2m2MA65hQhJef9CvIlLBKstp58boH07Uk1jRs1tYCTw2CAdAif
zrEU7tkPtlUY7z1aPz54AhAPkykiK5exDuEMj4EEF6ZRDdezNAzq84c5AquQX+ru
5dTbSxw2xnd5L0c+nd3yhI1uXTY/w7qgxj6Mnml/U/0m8ZWSu4loNcuSeAZpOx5T
8JXx5Y9DplpnVkOFq9pSchPgIftHQyeTuMsCQHmbjBfEKglzNRy9ZS/RzGsXw4Pt
9pCPynMgOodA5XQ7tOgMbmnWXxkwFuYCmnjsjRjSJnSPj5AMqIELQ9Mh2HDQnvKM
04AM1Rw8z8Y+LYTde1waJqkyFrhYQ36sLSl2UMzLolUdV/9iOwLL/IqKfVrKwUjx
otlwcsZ10OsZ915M3mWjkt+lNcrhC3lROiHxbT7kT+rWhf7o+iquLxamMAkFYIfd
OcD3bpPuAibE063FpW5cEJGQ3op9dfKmtL/XBQZVKxFtgvTEkGliDDj0q//aQFyV
TtFbYGnTPoeHezukjGn1uAqkQ/ZOTMLMlj1oUH2o9UqvyWjcFYB+eMsQo67BLqkE
Jz1fgTs8AOf0nZE5nzApugLKtoTEo1i2ZqX74ZIpNcC749+hpRHBWkE+HjHY4A0d
vBknBpW+NXkBaX3nMEdc6bJ5YD9mKTQJc0qIbrawSsPjmwGYMMJmrDlUgjtAKaun
yJDe5toXa2KWQ3zsYsIF/T2TwL+iBC7nXiG0vJnPKvrqbv/wHqz2ETxLSvmwp+kX
0j8uBEkO67SdXT9Qq/M/VBhMnH01mU3MBfXnMIcWyeF9y2zVcFf2e2c6b0LvhWuZ
shxrhkBl7oEEuHFVxB3RR6eo1ucv++sPxWfBK9HGkS3Mt9lY/XG6YSYRfSzq92Uo
SQcoeTssZNNtGGfB8NuFkO52HB+zqxZu9ranQK7tBk3fjp6i7Zkmm3/GlkunyPWL
6sCQwJMwvi+qZMTRuEEFUPYpMhwaYBDUBppd5GVdMJ2ne29i8oyvvHC5qT2VR9GG
Q7BVoI8+p/z6o7RAVIWAj+1PkARFvrgNqksSc7jT7Ikpx/A3Oi46uB//3uZlw/6i
rR+QEw6TenhG/5czMuHCHIq671WWeZUCWHkaGg97s8m4n0NIySCKhfkzfSPSBjBR
/jjN8l8K5vNMotuUXOwg0Gc3mkZi79bTNWRIuRy0Wf7KENp4edpJJh5p3wLF9QhL
kU14thVkaRJpR8VvMsNEdokfjt9efpNr2GVGCVdf7lfi4CvUWpnI8dGQO0u76wC9
Gt1RyRwCJVCN4dJgVZeWAR/sU8j19whgZSc2v6KIvjbHZm3NuUh07yZkzLYyhIm4
y+4MsjCmycGPeZcW0jV85S6/Ph0/dpZqNxyfhlL3cU0/thMY4SWuxzGaZdPn74U9
d6m4w01MY6T1H7CvQclfnz9WKTjxVI/SsSRta0in1MpygyPOgmxb1trx2rCjy4Jg
keEYh2EW+tTnJxYAfGioUuwOD7t9XZV9K9TPzPF8o+tHdqMQFTD1TrjWthmwUlxj
yEQmmGr70Uffn4ai/5cDQ1az/Vuv8iuYgaq/Uurtpewb6aRh4GR8Or+Q/BDDaUtM
svRXES90uK+/xTqFEp8xCtwdnuDbt/+Ud6e6reWl3iTmuqtoD+T12EdBMRN/Gisg
98cJc+hcC9dVd3tV+73Ewv9FmfEBJAcD/nMmrqvwXWEwgV1LxmoB527anhCdQDt2
tDZxLK/BPFxsjW7m1SEu4RV+23+t800nOIODsArgQ33QMLvZPBISnve8U/A9XlNM
wAWGBfRsRUTFDmRbByZIXmZPm0axVWBDKY6u8LPPyDHjOIYT/ZQpxcDlh3kzrYDe
WoyfwChnzHWcwpZMZDEBan/Zb5JGKFJ7PNq2BzQbK0KHuZSthL8hVE7LSjxm40or
VfGzphBxrE4VoDQ1Nf8nfyvXvx5aOuGO2TzpZ+/o7hsrqOmCZxlqnXG4MsEKgNMt
8H+wwJ8nHYNLLb1b9hFyMrIT+ihTuoWXWpgXt44jodKcIokEOfdkWK2Jymo7KKAT
BCOY9A6tqJkPWwvIA/wE/bTSJKoWF5J2UbRLO4uJJKstUbMgqjLpNQjM2jRABVYX
hLNvef3hSLkbPL5+fszWKCLhfL+rf3ZImIdxWJkbQf//rFT8BYsOZoFAqde6NAON
IHnxFY/aQI04doAVx/x4QFyeTIeA2EK2/At/uvPtf0Ffjm7PTPLf/PRSwbnYZ7x6
ASjgD563Me9RDc43nBgLx3qkso+hxGovwQgkbZFo2xWAxNxgQPBkZJtDYlerVe+V
HDPV1qoBcQJNnDKXghU8fBf9AYRa4mfazyzaC6D5BP70KZHCInlluiqMqmz9NW/E
zsZb1zkI4fVzxzhS14NnhIIoTz90FfYiax/lbABEKqbQ8p/QfSDyVryoRXhpnhcZ
JOAaBvy60gHiwFUKpGU7ex5WEV0zzsnw76HXlJuSkLT9UWwvEwoglUon1djT2U16
RAu5/HbS6Mvut56kZ+fKxsNM6gk8cqIxEZKqhaMahVtmyURk+Qb8O34mTOh2WVSM
crj2AePC3ULeTds/ov5zlMimI2Y6jg5aB7iZAqsLssZd+x0KMvI0rRgmBc3a/gRy
VoLPHQ8Pzjod/TEOlaYkCsLWAjJamPtNZixNEw0j9yF6pPxFv6IW71v4QygYZUww
7ETYdjiZUUKaNxNvh4akxYATpCzW3s7zNANeBjZoPIDOCIT0Of41YrfL26GSLtuO
Vx80rWk3XGcLmpOjWIqxeFTf6AsIetJUSPkrjeuLTe0JlYe9hFSpUZJ16bPSotv9
1oS2//nSu5qHEESL/YbrozSgXdc0LSxrd5n+BrwaX1hwj6L+8I2NqpsOMrY20gL3
Ij+X6B+eQWUioG8RluVagHuL5F5JbwSZFww0bIORHEoiSuBsbZDWAFUg+job4RAh
Ffpmb5387zZ3Lp1dfRtzCh6+kmAHchUOrMZlj0EUZp46cIIm6CfwzkF7BvcosrNR
UsdSDeHe1LYKL4lO30Pt0B9AkvqOIeFwaGAzdPClhHn8dVEiPzT3iQRVpjkq6X4F
h/JmTLzoWxzOC5VJt+G1C6ZdZgBOAWHC9MyRZEl/jTnCvKNTjLgm4hTuPBK3WyFl
WG64CagvJlBcMxNtWx9QhgyD/8GPKuBv6z5otjJ2QLAyIXzh8UT1p0JHo4Oz70Oe
00mD6Uv+GPhNx+mo/u+jy23N6Mtw69uv4aAb4bNBwUzq09tvL5U2TyUIp5JzYxET
0oJjI8NKxc4Wec8tvjdGc+wuIKtRj61yUGG+jKpDTt7dIRZAvIvoKrvdszLU3J+Z
b9p4x1fq4npWLcyID5Cq9Fu2RliM1eA05RkcOLROy9YpOXnDkmqui/3VRbN7B4xC
uc9wQ+tvzLfSHenW5OB7IseC0HpwfkZ7y64PqpY8b1RMRmZM2T4G8W90d02AWeka
+W4jM9o8gkDiTj9o1utpRxO3Koqi70ZiHuqCLaZXtWROX0ebhgrFFF6vO9dGKuKu
22LctQJBtH9VTgfOdf8+UmsdJfNLf4PqzKir/m5ruwfQ0dCWe0f4C7eM224Keni+
z8uLBYucPrUsjC9dC6mB2zI5JGSiWYpEXks50gVAZEMVc7NYuoqmeAepp63QToQO
ifhrmT1d1c3BMXSlxZYB7her8VAIwCXuypGRkFW0J397S+YjpLKioWZzarqeaBVB
FRUeS4JSCJDyuVgX7iiH/203AHwoAVAw+zPfwxYBBcBCJEq1arXiTUZhouPYWXOf
Pn/iOFHdc/Opb1mfOfA/YktANvUpML5QWBPZiEFnb7bl8cn+YmVmIBrCC/9Usv25
BWf/qGn6k70dq3pFVxpkC9Ik0J9Hlj58NBTxrPTnK3prJ6wN5PN7u082kyH0MgVI
z7Mx8UDonLx6Mw+sodOop4txp/kxxrdRkUmxlbtsMdcFZ049jaymR01r9OMkWp3C
jAd0Of6EkTtTRoKHuUYjsgObG0ttzKlLwNMSws0Y+I9XFyZehc0WVqkEXAw6Z+ix
o1LV6bECGjP0J2cR94je7l8ZwHP1jcAa2WYudeWUR6Wtdxg5SZgsM9XsRxdGLkrV
X9xtoOn8t9d6Dee33qlHvQZMi4HeTD3XZvhBL6sDObKz0Y8ji+Cap7o8aniMeeeV
EiywzF7cwpjemHChSOSHLtNPZJHXnMwIjAFEGo7oT0RjX3308exqY0FFDR3cFHj2
Toggf+Cx3Ab9DjncmVPxRklPoDyAgZ0/ZcBcugeq0CxvRGsOsXhabP/4O7ufhBoE
RPITa2EpnFr6Q9RvMS5OwWaSIxzldDg5ShKekXeZx4u033yFpwQp3Xg/PE+f7V/v
vydMlcvrer/i2QUIiBxWtxwMInXzAWF5W2re/bgzVG7RNYTy8W2KZpdnbR5fEX6A
Pt1s/k5kGg5KarUVqKeaUXOawBzgnKfdkLqpnPhmVhDpMKTt86Fz12sZxkmFLSwl
5uTsnAO3W6Pk1NupUS5Ydi4rdAfZDt5eSj9NN57gWsGmSYReIDoSX82sdeVPOLhW
8++C3OP8gmKQ9IzcSKkiMzk7N47V4yfZwUMW9WZcZGkXEq3K5pVBinW9slQuZQfj
M5Thigu1S65lnltJR+tbdsxTyC9nb0JmeB+GSOMmeB3E2XpI+Ubz/3gKTe+Ydsmz
o9156z03MHE3qUdKBDOioZYOTj1JH6fOH23zzy913xt86l+w6uJPQYPnk7rBH22e
w3Do8fuvvbZL3P1cje/Z6ynTR3e7rsXZ/eDpUWXKC0j7CAw/VulyubCXr+Q6JXti
gLcJEn/JhPpBHpP67WgM/oBiGjAyr/zgobtaTtzxcSs5FvelE1UsdAzYK13+wghL
BTJyRIL8fjrbaHKBoShvRnkRqVw7hmUZBt0BnGLwGiAZ1NSi83RPs4z7x3dBwT1y
a4hyq13y9MnLjX8c3xhLVzhzm0hPr0vyp28LrJZf5JBLLpnStVU3B1JKOuiAK9Og
lRA1eXeb3MoJmQrBiojhH44gAKSqJeW+MsLieXEf/HeOTZchN0Nmr754q7qeDFve
WQjrfTzNeDeG/3JQVVvRZMqo7HwoVLlHjcONPr/1/KTTIaoErc2VEBRoMAWM8ecf
m4PuyYHGQCZ3qwivt6cX+RcU/YCUbzxz82tNS2JfJ8Eyip5gTFUiITm0mCHL1UfL
VQajvu5qd0uCXqLw8hOGpaeza25tHJsm/Y+BWxpkxVQUC/Ti3cUcqBf4bhac9U5X
uP7WtNsff0AkZXSp7g3W+Z6uIF10tGHIwzjLhqoJA6A23zQaFRCRL6kpsKBOlUSP
hH3VmHqMfMBXZzjfI5Xlujqj+Q+yb+IAQ9YMBqUCJHhoN64x9FMMZa1ZtfOIddQt
85ZHQYT9amC3qh/eJMYg/SgOEvk7KY05AxKhMWT3zdvFVBoKA5s7AoC5zQ3QIwvc
Os+/Hum0qS2WQjzBe8ILE48wY8ONA+sTDby6FypahgO4b79VVAidvl8rro9aUa5a
G7bkGdc3j/bkr/xCxEjhavv8Y0P7r8lBMeZaqF82DUbGrNVmXqnMQG/nnj4bAZDU
nt5OOVuw7AMVmak2LQWXsbMP0kYrfnQ3A1SdL1k9APJxH0isyZ/8tBb3QkAZKdf9
6bnddBI8VOoZoenEKgI7agRLYMkRmDgn2DLTcjJPpQvKygr/CalC2dXFDh5lwU46
EXAHt5ntjijI/UoMmZ/yNopcwmiFRtJ6CXYTTAz6KNQRTyakJPdusCiBRFyR3BE2
CaMUcv0NxpcA3T3v4SErK0OovpeJUEjlt6ZNIZ7+l3Bgvij0OHrlZAtvtqmaRZ1r
ofd7A9FSylWZvX/CzU87xXjY65PvxYfbaRL0UQ/Iz9DTTj+1IUYT3uqRr52FlMIT
C9D9J62v//GXXh7jY7+Yfo4RUv6hXm5H2hbmqMI5QeK41yIGtuKpJjY0aJAVc+eK
XYsInlpCtnsDkwUvABqo0m8zPhHvwBQ0981u3pSblv1TYjKH5xJGzDkNo1VT6DtY
IQ1F5ASAVAKYXk+X3hfZabir3cypX8qGnlCbY7C0YA+6uHGKfyGBqZ2kAj2GFggL
UQiNh6GhxVhAyBUi6jF7h5Lc2nlGlOipQbh05BcVw07cbuDRcyeMjQTw22fPKTEx
u9vMzEO5bSAWIYAcdJq2RXYdcFhN591cl+1byzLrlW3OaDQH+gJefn4cI6nbpBjJ
PAUf7DpvZsWRea0XLeUckrNfw/2PT3a0GvldS5WL48S8q5iy39EYYwZkucG4ghCC
JfelELjCU8qdbcqvvXpXQh3mJb0gveflQRZvw7Q6tBu0rJabuF25LtCWWb9If8kO
pwybQrV14jj5jLWODOv5mzgHDYmReXZGT5UFG1sOev2DdRKLzh1ff0H5FrFIWFra
04mhbJxhja+dhEizUb10CniQczFdvcIFyYL/Y1MTqX+UscvZAuk1VUHOfIez49jY
GxVYlp5f8JK6rTlYeY+WgZfYbkGr73uhZtMrR/+whm8WDOAhE8SqP14/bos52FQo
6Q3RXxlQOpWC54AFaFQPuF7JCe0clNG96syR0nGnu+DVoqCxPAD2a0w+KkHI6yr7
Dx4TSzdtWBjxjtVLsX4XLm0OicoGNASD8//TeGOOIpZW9RV0A3mShd3KHBUMqSfP
PIUlUHvMAoonU189K0+01PbYXVwacr2M34CE4+uF3jvqOBpIqf1NmywB1rWgm2kA
Xkdk2Yje9rPamY3y437a6x5YUokTadeik1+yDTiTURuSGrDAfGeLRB1V6tWITxKY
Vnu+0exwJP29SwUfXaJpcjaL5dZeEj8ZZzzbDS7PBQMeNADVaxc/tpQOydSI+SLa
djlwCLFKysrZcKbkBrN7YgmXKi+gq/NdBLT8eWpdJOHkQrg9ACE8ToaWtIfvHPDh
VhxL/cFF5XtZDS1KtiQlNgYfN9ccZb9/CF58kUpjtmo1ZNrM48RidpqieIqb6d3P
Y4+aeUueSPM7BgVb5R3JLN6EJi7LpgbntRZX6CzP23TO/XXjt7luiIWZZzyXiuys
u9+QkFShjnozR60uQNThSOwMYAZf+IfzeQVmp5Wzr763kZAFBZF/HTrY2Fw37D67
lLrR8sEUQvos4EOsmwMFvKcuXAOgV6OPgKtJdz7N8s3NGg3h/4VzoSyKCtacotaj
8WXFim6J18P1RTB7NKFAgJHL9hgpLZBbwFw+3CocCJqWNNmRxANQAizIMXVaXI7u
WvJkfRSBbrouuOegZ2pV4TMYA0hUnTMFWk+TAhiEN0OsRo+W6PIaxZxDQR+r3ZRO
xTHGXJRuWibC/NuEZJQfEMqVRhKt2EJRy/hS/xeZDK9/pRjIZ1YvY850k3Ai0ceC
ylu2MmaMR3opfKEZZnfULNt6XOvbe7sAi/8RnnDnh+aQ2zsAAdDC0SG0uqEYymZ5
btVeoexfa7glykhz8hKCbO3WS1AJrDkg7gYA5uzq/GeuI98q0ypgyh4acQpfDNcX
gh1kSxUnp7fhTQGUZwx8fuvWK75erXzNl4jF08J9xNPCoeZjYAWRCGdwYMAyvrWz
+eD0K7IKu0S585XXtrsDI/wAFy1ti6RuE0RHqfe9fW9kTIljf03ZRvOmiWCAjGsi
GsQYm7Y07zZqH8KR/Gb1wic666erC1HKHpDweidl8f+vynHD8WORnfcTXmACfDBZ
IxfpQcAb7FoY1aCp7Eo8jngb522kG2yPJnKPzZHDuzDw5E+u7irlDP9eQSraANuA
9hwx6bufXHBjWj18e67MaBy7eAPzCbkBqjYzSVz1Eq/ukGLEzYTaIiYbDp3VbghZ
aNdR7F3XrBtQSKqz5p1kQykk7jJhGpAdQPKC0uz4QsFsefL0W3yy+Yy3ohpjwcDa
gNoANpLSeI081dyzfYnIdDUmEYlSbGbyqkUPVVfp76SLR6/GBNsvKAV4ywjJ1Ofk
UNOGP7wCkHvk4TAdIAWOr1tNKocRStuhNGClSny4f8N/aXA6jK9RKKCGuJg73CT0
ifG/cfG5ILKy/sRIVCLVP1juwy8M6j7TtaRxxRYGE3gZ3I2p4vU7cOKFkz+9C92o
YOLWKc0Huwg5XtWtpsP9efC8cSTWS8D319J9UW/SYX9kHa+8oAzOA8WgLA7zItKL
D7sklNbRP9hTITk/65UkaeU00XptJHe6yUaA5+RTiPVWlSx48DQvHuMKK/T3dLMR
YaWz2ExvyzjddkG3YOtKQeQl4QFhN8ZF0FaDtVlbNVrsgSDP7anPvDn6GpSmHxwL
zHttqfscO8yR1flC92COxGZ+lc/nZXHFEwCEkyovYpsoLPb1qXX+TKIVxGCyLGao
dBJ7qR4E3+N5gtL+6KtiUj0wxbabwyR0IWG0x2rLMcT1FafW3sNk+MicVQmO7+Tf
5JzobwHUvq6S/+JC7g/z0diCjm8kQju2dV7tcD7w4EY9dnY/blpSozJ0TV7+XrWJ
5HyrU2mojwMcb0qrsIX2eOQm4bom7SvodCyF+fMoi5V9SkAsWVO/aKZrbLqDviIn
r1mUKcg5HwR+DSNl7dybb1t3P9PNJ4LiIAd/YuYVNueKVM/opGQuw5G4JZla3Ijv
22eBwu9gQ/+BIY+nZ2sHLTWVjle5kRIuZqzf3naZP5Brx0nfDoiT0LuQBrawGSgO
Cb1gjG5a0aGHCExMlQzlqM/pEVUFID+mT5SOo/hksptJ4a29nKlfg0mRWZWZgxts
/HVLd6nWJxTVIRqQCQeasrXam1bdvn4jmykF4YyeDYY+kuXppTTZlhCsHqkt15Me
0hp/Qwkv98rjMZ670lazpZ9aUwsJ+9osA7J/oNEEJzxm2u/CZVQHa+V9Ixy72Dz2
RtXjYaI2MTGtWs6ugI/it7fgJVQ0xZzPE9UAddVofbfjbalH3w4I7xRFeXDxLwas
Ppfsie88vkgHJNXEG8ZuDGSw1Z5X0/gBKOYRCKU95DetWc5epbQRboMl/d//BJDl
2RNfkLesF+4Jszf67QVwngXON4uVcoNyKfGR5Fr3s/z2RezM+pQpqsE4qiwiWpBS
PSuWKVj9dFhu3A60cSGLO/zjPSYDtGvZQDKLvsV5/rH+UL9EL3BMhTUKADRvt9dC
oxoJpjSfiaMTuOGzo7EieJ3sUZxSUfPplYhAEVoAVoknV9UYAcrHWFubkDrkDOPg
7XBGSsxT5aSQNVIAF/bTtd96J8WhiEI9D3mFxCIAIswqMdHkydhcJCMMdCIwq4gJ
t6eOMKqebMDc3hpmTZTRwTGWj//jETl79blz2Yoq5ABTp3ZV3O7dd2sTshlFvRmp
OrcvL/tSBmtMAu86fIhCXr5EjEbwPRBEue3jqr588FMc64X13XIbv3tBMTie7okQ
pS+BbdI8lXCKsJ75IomkyBGs0AnWa69rrgHQc8qy9XQq1VNIDIT+LQjzqCYRaDj0
JOE715kI1JJs6QXJ4/gSRfc/qdC/LN/i/k8TZrMQMISnwoGn4qWWPDp3ekNqTd4K
GNND2SNA3uAdCvyv76fWYZlO6tOBLPiqLzdXKoU1O3NTQQauSywzNwrldBZm+GZE
U2GPw1yvFs6dnp3fpn0UhoHJAcgo3d+y2fDdtYfc2JVCCPEoHvw6XC4VIqFStEbB
kI4gXXh1TrghFg3Ox59pEd/6tufqUllLC3/4ae+Asury/ehOiWClGC2oTPGr/280
8IjbAjTNqC5u7m4X/DBNsURglYDuDBgRLwz+79V/XYWxqRRdyFTzPc6+0KVojqnn
HXYnWzVYuAK6yIyXzbyo4lu8Q2lTAfBrCJ/CTuWU72uv/JoNvwc01Iq5RzS/hu9Z
Km0l2rLNQvkMJ6aLHnshVloz6vPzsYhFWtejszWrQgC9c/yXp2sVhq5Yw3P6oili
bezz/F5wsQJkT5lB5dCjVQ4gKBN+GhDWP5R0teFEZSgsTYSFY4uvzFNRGyDKRv0u
fjNl3B/nOPvh7hGqxSkTfZ/CmkKrtF5DUcqBj+NT8DXPqcG9A32FJRORBsJJ79tI
OuwE8hDaqUMY+DfFCTZ4dZjS2pSbcwiO3X03Bo0Ufz1z6pksFldMIsx9lkrKWx0i
TsiGp3QZAdvdMaOIgY9B/FSlT5wb+bngUiY/g6p2mfq6yU+zzd7L9cle8go3u1b0
4iqVcgCb7IZAl4Z+P+7K53ACKfs02AZAQzdXBPfHbd6qA6oboDywrR6pdIex4umc
JOTC92fcbUSXQgkUT5+PCX0baT/hTxGelxez0LKUeZbb8L+J0dDGcjY8ONEng/wg
erg2iZ+3VZRIOxLhzL5UPQRZqX17/eP4QXRj7Mh6hEU89jmw7u6NxkQeRM8QTbpd
hyueCes0HZwjDDRf7xpHvJYCiFoMwJiSwluqPjgBg4+vDJuafsKckeEJsEC4t3Um
Rtg6U7rzosgNnacMm6Frzg+W+CU7V8Ni2s2xgwR8GInwRLE7BC4s47QuldbH500+
gqrdPVlEZJc+Tdb2+6D4XoSv6ofmjV4TvTpceOLEKWjnZokQMnwG068rJaOWZDY2
eyVOshh3djWEMA2MWYoisowR7x5pzUGLZv5y4nm67mlBP1tLiEB8qs0uR14853eo
XqAKnAcWe1qUWyM1A6o5tXDpWepx1ImwtCMDScjDszeNCfoAoZEbNIvoFYldN4rm
B0B8nm7CU6f2htVgQWYK8kcmkkMLD7oPeBU5ke779IyXKhjasmO2KlW7wnMO3tgc
R0Z2UHNTE8qqS3xpe4iZTSHtopZaBZ9SzrA3GEsVumMkh4m0UPXezkbyeRB/KH+t
4FsKsrai7HYFcUYQfhEy0fh0ehtvNb+v8F8owig3a+LCekZdjGvCENC2PoPDlN27
HNr9PsI9Q0WbhkeCZubiElxs8/IWVb8GrX6FbzjeQRHeEb0TSfCMyqGvZtIZBXU3
4oLZWh97VAJf7i6Byjfue+6sUmryxNt2NDxkvgtjIGzeHftzb+UPlETESJkXEm6d
TAPmCxr7EgRGUOB0epOXXkBBgJBxPMRQqYM2K8lLLVhC5VygVb6le/pgDgHD0sMr
JYIF5o7Bf2T0dPOfm0jBmQW30tzhSMx+Vx8ZnNbxMbW7zp9Ycri3qvFu6Ppf2Xfx
QddzpOmWlZkz7QQ8J5Bhdr1dFo9VGcfKt8L/A4tnRCratHcVMRVSQbvkG+zdSYIJ
+pZ6NflBQlzqm0B/BCQUgcZAn1WgFrdJHFRdNSOviYfhpBnsE0br79Nf8kQr14+O
PYV8DwiHCCN5b4SpbzThS3N/xiMqMpGFzYAtW/b7D0F5mkihTrp1IbprNg2Z5xJz
i5pB9VUdAou+qnED1pGvAd9VDpvMErqD1iOlUXxHkN2mpu9IGyjOckKOrbAV78dP
lm7uVK9erpKItaVPZKssZHJklYOK6TpWHvfWgng+2/5a5v6UbPWZE35rGhq12gQ1
7XQ4XfjyQJ/sofkJLzfP2fcnEVTYIvdMS9/PmSRev5dk3GOJ9++lOBnaq6sTrRFj
nCzxn6pRfn718rm4/4uutQkLIjHF+B/xC/tvg1/dAsUaFAUyAJZ9OlMxKuvZdeQa
VugeEyiwjOZqCdmQ9AKz3hlnNBNaSDt9hvzujjFGa/qgxVuzgZoZD1TSycBreCOI
hKkVN5MqTwOeDaRtVgXwJye3WcNG5ELcn5fusNoTS//gEZwFKGlGaX+l8bIs7Mie
bd61mOG1eh8mqyMuIUk4hPp0+l5Q5AKd2OYLviuCeQlVbL2WEbcTcIzVk+OXcLoQ
DcsVF4EUgTIPKqzty76CRO4kk1uGfcDDbmkOZWG9Y9igx8Bs2mdYWhPkP1xRtCxW
FWFxm6C9DNmwYXC7AWyXsN6vnI8XxbZ+tjGbP/o4m8rNY+GUoK7ZtGhq29jdr4kv
ildtu1HEldB2aDt0AOTlKn6jwb0L/xoav6/5jMR9WF9LPcPu6r35hlw1pwWjaEAO
YnV0ynqMleEwQE68uK3xiDqmcKK4KztOXSDWJFpLm5UnRoyXcm4ZkBy8rSd4Jkwn
yDzeeWOvQ6HcJoMen6+EkmJPsnPwyfsjSwmAsGyqeqx7uXNK1xJ4lV3Pqj4jwWQF
Tm/BUbYvU0aL2ct3HJJ1zfWEmDvRETWKAcYqV8A5iQFjnnzAdnepQwyo4heNAaX1
oyI/tsMMQwqOJSjV6L6iatxCcCYccY4ZWJyfFftl+3Qxw5q/yRaPOeC67lTK15Ch
rddw7uP0PVwFdZo3/iUOnQV6r6xpk4gx1DA0Bf15L/4ImqYWxdWCUibhg155ZKtP
60A7x3qG7E7WewNIxvsVaYH+ZYgpvBVOp4EVuWsanrUBkVVpf4OWaRwSf3gy8XZ8
b0SY8IHZpG2PAC0/pTwrS/GQq0xO+zgBzjpelkMN4bI+Mw0KusiMOLf2ujdi3IxY
ONRug6tTr52U42PT4PLStwVXY+CMGVtMAkslcLcx+m1o3/ANiOAuSBt4AsS+r//K
dO2GVI0cNq0Dgmcia+cgwiZYJWQTxHC4HAXOv2apNcJjQo0LAhN6WZfYvs+8X2mm
NSSf+FHtOCWUjgkii84tF8Jro+El53JAvQRj4EAw2UOQlBeP+X1tc6n7ufzepXtJ
4ljcCARDbn8S1nqdwQ/M8d0ce+UCSWgkqQ9j5co8HR3cmkLaLYAfP1R9DWN5ZeC+
KqvJXeSIz/z9902f32nMIlLP1K/L0TJywqdj2wWNEROKYeFgCwpxlUKWLHFrTBCT
mlOFQEIAsAemvPqwVAEAebRF4agiaBsjayhgkwVey/m83pqPC08yzOwJ2CIi0BM/
5SMUmZXJ3D0HwuTRCM3Tu1wD346ZnbD+rALloAbTnlYFligeD2nNYh+NNEAifylQ
s3TpDDo3Ftyb7rRDYwn15ellORbTi8w4StPDrKKFmPEQY7YubAPpqKnpgA7x9a/H
7oAibtxhX0OHMgUys0TgoziHf2y1qGQ3YMArkJBsNBBErUieIs1/Kk/yWaf3ShwP
chNhOHTVqlJLqYapzu/vdinau3mg9bPCKECJku1+5opRVZ5rcAwEuOKJN0ieC/7p
xpVGh1Zd4sbaAoK9WDMvr0EDCDMsubtcdvT9rsTnB97/8ZA4R+bFM+MIxYSiVi9A
KDXXmArKLjHhXu5NIywUYrD/l0h89yp4ydx0jrKCvPaiV/lVbWZq89aNE3nuYTVk
fnDMfpaAcvYLIAfOxm7WDfNv8Y/l+kehSlSTgSANFEwtnoHLKaV8XbZq/gMCJ+Uj
VJmfh22zODaWyyUs0uvo2rUBn2JG8jX8gEqGWUWUrtDwJqLIFDxeIEuEm4txzynQ
DukC/YbYzotx4POvQ3BdlTMhCG18yPLc7CZc+9g1iEMoMz5g+59vxDDcDpx2pGqq
O5digpvr5/UhEfFB8zQa2jrFp8rt6eLAc/6tSUal4G735d+KAFq+/yizzRZuty7M
3ITeZaR7zimxrRuRfnq1/cfYVNxPVb66jHpQ3y6/9WIezzdHw2hOhnndIXbYgwS1
nyu+PTB9QXAnu76StE8BHg/cnUYXaS6UvRGjjvBl33XhD1AeaaYzlHO4mMY1taKU
ZgKqci2xNYBD3QUTB7OXRejHiJAJLFN1I9uldtN3VthBP9tPIXMECQmafCWPPamH
Ev+Ey+LsPTRcpP4WJ7ETwJ49CLbOClHsjBH+nSctZVXAJ4xi36K6WEIuGEL8fMdd
Aam36wszb3FUuCiNJR81ETsT5GZrifmD76Thk1ScL0mC8wfVN4OydS0kFzQ27sPW
PbYcSUTd889P+KcL2sUaZ1MglEdbRlmYAXd+st415PJylFdQJkzez2DDj32xrQcs
wR4twsCnXvnj2ilknY8LA5SeEadgiNpDn6i+wYLAIxAbb1CsIjrjhSYmIkrT+p2l
aL/6RRJShT0UwEb+8rzzrzmn9P5HqJYQmIp7l3zKnvqnIxLxziVE3uJAVNtFcaGB
dfIHx5gt173tv9HBE77KHHomEB0tAx9XYgS8FmYl76LYqYx2JMWhE8qgUaOXoeAU
GZ5j4Z0IIgHTP/TfM7sBw7bFF9NTF1h7xpepyOaX4L1ZCt2nCJAEKfI44zzrVfo7
GC8bZ6/8JiIseJHIDQyKVpizv1WxdbuYxKZNe2O3L/VFM/qfOmUOabXSv6JfvcMp
kD1/Ag9vQh9qLh0MBGYm77rJJEUFlqrrZSTDK75syoYLfoxOe7G0NuazCiVflH1f
l4xjUggGZZGUDWOUrHLTRiKEi5A26lRNCVRjWA1eWJixxeY66TlshK9uao/21WjQ
0pLYPFYmZSvODlyRhdYX2sy1c4YzhOqw1NNuGLdmAht9tiw5QD83UPFR1dfRXeI2
skSFTmiNz5a+AwMydp76BoCObl1pF3FQplV/F/WuR8IEybj0S87WUmgC4mfceYnH
sjTbdZgzxCijLuV4BQsIN1ByWqFX5womaFjV0CpxFHc483gMlGTL7iD5VeKKQQ65
2/iDlQsHeDoQAzVJSZaiESDlHU/776Vjo6CS4dmE3VvkUdccX8FpPfD2f/qZJeTD
ncrzjXv8G6F07O1G6aA2HADR/HkVobZS4YjCLTeBsASPbUsHT5YZsuL4te4qM3Ww
pM5XL5KTK9wKkSUTh7/JvZdIsAMs0iBcy61t81yz9LIrdr7tPlw3OVhKHkVw5Eag
Lo+oGOj8t1QLmF/jfJz34wEa0yjwZDEDARM3v7v78mFFiTs+1pz9qPtpq7gLKelA
6xBORcjAYbP3ZeB2agkWrd89+I6naB+Ym20mZr5WIjaXzEpqK6soGbcnM/aJKjwh
TWZvU+PjDzWC6vO5+4MwZdunLo+PtQ09ZKcirPfctnclJqjWsDmatDV9BxzainMP
zxUpQT77ZpUY8/kQ14NyaC3DtdO52zrqX6573jE9WuTFpLnO5ksA6x4UwNIO26bv
s+YPLrixgvGEZyXKAeEmd6DsAkEFZDfZZkeqMBlnMVY65n8qPgYqEGj2VudXcgYG
jDOFana1JVpMWYkZ8hQLk4V/yhYmX+10Pm5VXxUCDZ3IjfNbF6cnWMcp+hH1ULdp
OC3ld/K7mxHoutP3w3CxeTNIAnF1/qbAJioYN42qSzAy7PYeOpo0WLLpQdCn69Oh
Ek7jv9nV9FYNbr7mBNnFdzGcsZIgjXs5EiIj6gOIb9bIfBzUkVWlSsOiW5JS2emb
VPUk6iWxTBsBNGxYL1iq6SwqVL5gQNb4Vo8GDsLN4VSSSHN2e+MbCeVMFw2Fo27J
heG4mP/iNHi0GunP4t88XPCnT+cRQFWY52VfygDRvmW/MhDehuQzYrrqZ7h5W41h
Hfs3PI7b5Vu31mICxOZZ/A1yu31c+Fet0/4PVvnj6aY7b4nBIzMXoQAbE8B3EpFk
ttfE1HGebHE8Tq7fQ0mPSSTJvLfb+sUbmT9KtSBlf/ntacoA1HiMA6Tl9XQA2WQG
yDHHe/l+cCnzFmfV6No1g7Uehx6WuR+hgeW0Ro2lhiCqS8oQQ4pbd2aLGwyTAurp
qzyV93OZVLQa6ejsq/tVILnP1QmwlTcxdtMcJI54WeOwvNhQwltM9Wx7lRX7ns1U
UE5WajfCdWbv+3dv60Th5cW2o5ZPdRpVyUUzh8+qJ24/2vJWpOcL0Sv7eEOpy4Rm
2w99HSzrO494s32ZMY8tli1aKnmcZ9KpHnp4qw3Y7r+83sICZAOrQ1il8r2uzkKn
/2Tc34BQmRi/TG1ZlKHG8/5qzWWEaSLBMl0TzUTL9U4yOcJ2tmgqZnDpgHZoTPBp
7iEegXwXd0hM1gH1XGCtGBIjBQ0I5HLhsAOeL3uTNUX7pk/SgqVIbwJ08XI2qILS
j3B5M3RLIkAFtiaHegFOm/QfIRHqonCs5kEofBeAEZvPkP0XBgJKOBsg/owPElkE
HgOZeSbJlty4Vyf3dXmalFx9XgERfHOxKZ+oqPBZlfriATwl8HNJFOKX9A/ypkWh
2cF00SE8a/dN0rscmrYIIm6EaZlT27UAVfwTiuOcjtthpt3pEgXbelpvAFYGeMpU
E5b/CA69J8vsqGiJtPT70tBRV7JoRf1jjsHLmgHdPG3pe4HuJXDestYLA0ST7mh/
BXD70Qva+n/Gbf0E6nhKEg78WWvynwQke8Q/nLFBzh2oOXXVGxyCiOtORSsQz3HK
heBaMgL2fTCM7LlrTiL5jjIzjn7WWlvrDreo0toun3qArnNtktwp/AYsncM/upNV
xcDsDyn5Gkw3YGqcGhKSVtGZS8g/EQgOcudtX0enP/IApMTf14p/d6hAU3iHsdwF
mjbpMlT2QkW0O1jauBKaTvj1rwZ/tNQI4lyD6x0nOomr8hKYdRhU4RLVgPnFpPmB
r4XgOIuU1equebFShodsz7DeIFLr/bmo2fVPhRbX4x8jhArIHZifYkhkssW+HkAe
AGk6XSLMksaJft21fjmuMW4sjb0+COov24viW49TFZSZLMxk0OsMWt+H6UWkI7dP
fVb2rbGA9nPhazZ0xbwmEoYaSScccnTU8x+9KAkcL6XEU4RlTbbia+pIPiyK5I3W
aDWYSiJ10hb5c3BBytiqSG997cudcCXcOe3YfDOTNyWv9ll3ivi+bHk+lW4X8ECU
BtlfAfZKTsmLyx9PhcuSVyAjGO3Uzr/F2M1TTDDCFJ9lKBGHhQOxlSfp7nejDCbx
53nkh7bMo3UJlb5oPd3iIKIGouyYJjXh4egcq0PZo8nL4uqq2Cw5z+a8irT0/mOr
JzGY6P0OXRra22T7ZtGWY6d/21XHRLAUlV44PtKexvSioqySwyDY1b1GQzqrOPJ6
6jUocj4YiNt7I3NTZgYWFEnz0hnB5tCyjysZ8RkW8/h1ZMqhmbSbX/S9VB6SxjrE
lDN7Oq+4PQIBmGwGtUspxWKP37fFeqLJzsL3t/7M3BGuyHsT6C/s1O6zmemwZQcm
GoZooMf5abJPUHyuKRp+hA67NKGLYfnXxZEnPulCYP8Zqn4X3HBUgM6gTy3F0o1D
hCEXpv3wXUiOsdKuBbw0qMxKLLhPfuDBuvyFKwLUmLW5dURemG00Pn9O/QUktLwd
rvkBvrqExY4heN4QOWGI/6jek6RZiKIqi/gli0nOoic1LPjq03u5jRXXtQZ49pkS
SLUWmKrNSQ39rCNHf2wn2Vn6pZhoGDX3l4mLOw6bhFwidDIMqCUgo9g+AsEeR2xE
OcNRGrxdws2uYfUvZtE1Bq4WAs+UgB9QFOSbgOa7suXLy0orxT5t9gmPoPxPK9vO
opcG3Q3ij7BJppBbyc5PI1Yk38Jx/Pqnb0qzWwFt+vSdYr1ugD5s+yvyzQ0Hq9Iq
jOmi161Pe29Cc/9amoRgupp7I1S472kqfonB6oFRsva/maWPxupm+KomDSGC/lMP
k4D1uJO8dC5ItQEMqcef7jHlglVC/n8kvmQJ0ox09Ime004vbxXcXY28oLp4egIZ
AIjd+fD1Bh7GauXQOtfrCXhg1e19RHpaw2IE0P1Ve+OzoiBar2JB5gbsJbASvZm2
PnqWQT2DTo3WVZ/qycKMnWGoIJnXMMo55WZOL08b1eu/93qEUmXZUNVwiHkBeKtw
bnArytmr1GIXQT1bfR32mbXs4rYPnxSUPyuzzO+HCfITEHPVg5sYF7LXUzlKt59J
ut+jWInz27+yoZkQDG19lComOp1YwLMcUMgni1ahgNDmNRrrUYLPtgDJU62xKoEt
2wU7OH3Xf/vqwZWxU9kYX4zhmdZWH6M8zAxy2gTfPae/3fnNTO+p/F5ij8NPhZhO
YCfPdgDP/1mYccvIGYD6aNxUgH5vw2vU2Dz/7oW4h2cIxe+cF2GI8OC29iUlSl2j
gktN20WMwoRbnmJHx/YcZM+61ZqqdSd0nlyUu7rMB+lfO+eE8k3rGANac3JK5VPZ
tgB+olVBEkNdjpTAs6IHNhmXuNEyScjvpl5eVjBg2slEjvw93SyDtiiJB0kPNcJP
/5h/zVpKzcmVHnzGWOuxYboNK+vqAJgS2owzO7TpiuATbDrEa4065/6/AiDJTxm9
ZQLPlM2x7YvPme5WbtqL5htKha1IAPo+NaVJf55tli0ocQQwGHcl1w6qvzFXCJ5q
WujqNINiqGeCzji47QNw4+CRjWbXITXEeaUJFjqmfxFoTwzII15+HnXmkaH/cq5d
IK6DXoQY72SqTtSr/LYQ27AmfnrcIFxMOdrj1j8AshiTL162JfnStqM02OUksAIL
OTUkNzZqM7GmUB9hhiJmT2L5dexyURJITLuoijiP08562WjrgPtrYEIgky9aE1FE
CAWnA6WH1Nc+3IbyeIGoynU1jY7gfzWNMIXDWclKdICLIOx0/MelOG37MZydCU8b
oQRFmF9ZQaYUq5F487bnymTKviyoFag53hz+S6vuqT3K8d0p1OP1sNg9DbaPC0G7
gOG7EFV2R3tDDxV7rVCnW6SldxE3RIghGL5OdUkwOl/EZue51/0KSWRylCnNDvRW
RMY63mWkpqDRoVfjXhSBb7G6FFpiQD63gtqU/b3/75hJPjtftbCbVoMjvEBFjy81
k0rxZibNzWCh5vEN92aHGBGzpPST0A5SPIu4zK5ycRLoMCXqq6xtnl36kKxH90cN
ClJje9f6l+iYZn3SNpwCqXAQhB5ffBteWJwxUM13vKGUKjPoDeSMiY/rnF2zc564
FaNuYqOwOK33iYJOcMDxaezyoSjsehoqQT1Nf/Bo8o/Q7S5W4HnQebhO3A8ITxd7
9PcLwf6Bsn1st86qIHgGE7cj+v218sRAD73XlvIVZs2/OnmZ1z7TeaZ3zXqiJAmV
Z4Tl9tZ/yPLTBa+aIuNVq75ejMFhCCm2DJkwZnOPisnWpNV8FEMZoX6S+W1giCB9
mwa08F2vwanhyQGfBU67VO9PDeRYemSjD3IGX2a0vhPE0GwoibKERh4O1d6kS+fk
PpCqBDvSbxH1EKipf1II3HBwMKyGqYfNoTaCYMZS310JPCRwPncN6o8fdivWMJTo
sWjuSFuWL/O5mTFdeInGZsTvlyWtabKYSpdz5DZ1vj8Tu1+QcCcbCpnVYylY5s6k
cgf1CRBL3OGawEucxN5Xfg8VZWPhUAyH25cCR/UPhuECWceAxa3FUJNPvQRj0Orr
kdzOFcHpRt05FN9lCky3i/Gr0+36yqwYrw/4vCrGPgsvWPsVun+FkKWmIV0pVWiJ
LnTgpX3f4CHLqFwJRK3gP2ZceLdHXotvuh4/Fx0FOkvtQGP27t3YZUnDBVMsUUPp
1zEeyh5bH0a2/wjOY8OU5XRMpuTur2dpWdiKHlCv6orFG0Aqfki+kmrZdB3VP5wk
c/A55S6Yw+yHbdnr44KQm1N7ZHXdETnZxuN5QW2drbsqViGC9tAdt042g+yik/oB
ze4mC/oWpPPkEW5pu1fC+4HcR40O5D755Knfa+BvA02QXSAFhfipXBzwv2lRawSp
CsWmuF45992bTnY1gvk/E690SU8KZbJudPK90NrQjGUJLBi9YSlb9sSI544EEk2K
iuWaL5f2oSUcJquhb/PRrWQO3OiXkiJF7cgQFQ2YWhiGYWQ7mSnV6DGgb348le5Z
xWY/KO7DursZtS/LNe036Iw+EmdeB1ILUMhk6JMjCeSQ+SL5eViBTh1iKUi+B6No
DM3mZnBtt83b5nwIe/E/slOAhBPAKOw2EK++bVt95WxIRVdWV6P5t1Hf1Z4jl7iW
3vk8JVZ72oBKZwN9EUoPDP0bo0mdA9Gv7iqKMkXBkVUuo8hVE7Rs5wdZUzY9+YrE
CGNB35umwLnoUrX8jzdbPegAVXgls/gRZQjxvJyMzLJtcnbuIgCm2gdxPic+dtzr
gpjs2fklu2CAa5FLI1ovrjPZ6CZ5wBbZohj+J/0qP4BQteprIv5Wt/2/eRLYQK/j
saYtE4iUNnHvVq3jWWkSJc/uctevetYwbks2Wf/S6PGdCGycRXfn38GrqwymJSZf
Qy6MBCcY2BYdIYVrAAmbfRemTOqLOxVW3Krdpzdd4ZYvQzdE5LuZBPYjVT7vnK57
7OQsF3Pr4FtJyibp8cFCsiG4c2JKn381DYiBU4FfX8vzzoaWHnJf7eEP3Rsk9HQx
lCTXgHLob7lUJhQY9XtPjySlhqEEju6+ZM9rdUFm5vyjCH+wD/+FarlooAuCwNR8
v9oHRl8n1BhU0QsTgIaqFrizCKpSOFqVb82RYM0qLth263p7/jvGucfvoiVCd1Qc
0kFCw4o3EW69OZPHjgPaHawxytFvmUfxXXXdbnhWEz24+AOBoWWoVRtOxowtuX+Z
fy64B4I7lnDWerurNKp1jaeCA7le6DE/EGJe03tvs8ES4bnj3FfVNA6CS7b/2XRh
xUmS8lGkAU7+fcSUbDVmxaYOmA3/1dva78GtzG6tMSrsm+Tk8ZklDnN+IlJoSjEB
fiaUASWhM5UKl9pi0n2BhXSCCbBaqaQL3KYk+zdW4XGoXn4FxM7ZJYR/cKhr3ykh
LTiZq+YE5Iplvwm2+gd1Xe+MQL7IWfaxaypZsnkDoYKM5TcgWM7XsqJ3yslIvTYZ
WD+gYounp/BjF7tQiWLOEIf/JiTtfB9PnnT1cvGT7hcqwSOxgBYBJA6DhaaZgRR4
y3lB0SAiGsiKrJlsq5EIrXbfrAo2fhWlflOSWVA23cskHHVB3AP5cwfs0GENt9Zd
nai1BJXiuUAxqRnHnh4q+8iPiCLdOvjXLCxN+R04TTfnzPeVkcfrxsfEi0TDTbmv
M6WoQhGwcvKNm8FWNcGeFs3zLfUI1ozcpVNEmqGxqT6X3TIjFrUC6uHugBNLuyp+
wgZkrl4FMLiTzIQiwP1JlE3KMfi2AyJP5yDFEYKPwvdEDPl6xKhX+3PM+Xlat2Ni
c0+LVvw71rdqsTbPYwcJBhRg+vU74HJIkqrjiiVOlI4KyQN8LLsZG3G3Y4uyF6oc
ALwvSLYqh6Te7tRERLm0yz91POZ1R1hdgc6/jgmcf4tY9vGWbIRPhAPxJofu3YoL
8futQCh8doyeA/e9ZtHiQUWpKFeu+0Xqtkgx4a2plvJCTVL/5Qiiukp6Bpr6viOg
D4drUIlR1MGLiiU8teJpYCFORht8UM2901TghgiNr3ckVAHoZan4RAXxbOmsBX9O
2Q3Puz8nF8GCFJ26HKKxfAPS/hRsMOiB0TiXh/XNnayXxymCbmlzkRSAJ9P22/b4
58s4vba4yNK7xt/qxJwGXzdGk64bhDoSMPNfE+F+zeqJbE5j7DfbyvzMil78gY3B
LbY9jdXEtrxfccXphOcetpaNDG3ZQgRD40N4E9n6CtZZ8K9CRGPV90r5XmAJQtWt
DzzkcegX5MqKCXmmkiyFOR/QjqY+9xzdoCEN7hkg6Y8irw9qYzTLcDWn2nzpBO/R
d42Rv6d6gtROCOMt+rb4XHXD/ckKRXGBl9MdRI0gvvteZsRBXsmfY0AXI/wH1CDS
GXWRYZeNnkBT3S5pYywPtlBMhFXyiDsDdmY38gi3y2htSboeqwDxOoLWI2q37ZZ8
m0ika3YWyZpovzmJTGdakF0mzYa+crl4JEq0GL060L7UIFVAY/emKIQ76Qqo0MUa
/WyYOdXRUdOTD0HFl1lgpOlNhL4K7z3isJL4EYjHVUcUjnMaIvtYhzTXz0Bcjpu4
6eOABiE9tXt///k5+1Mqs4lgIkhi11su1MPWEk96pKfw67VcpjLnZEf3F5uytDZY
Nz2cK0XMonO50xTFBDNYi3hqTl1prD/Cx+LKBsgjCnmBZjVoNQzQqS1/dft05+U2
oGK6wOenG1M9q+48QE59Pu/Fx8UklhvAEECGq2LAbfD3pCxi6NhF4XyrLClbqPni
6iPVIR4AssK69XeMLvl1mz3Yf6OOn126oKM0Oyi7KQDgG/Q5YZS1D6OEmYg0lRZi
xhjhZs6vnnsagW1zpFi/jzrmluvV4qOgj3+Qnl25r+adLEvzZEokyXI+3+uJruyZ
U0rrx1KL9aw0FMKBxJw8WmJxaHcx9NOd2eDG1GsLjpiZY950qxAr6ayKjgUm1pek
JbBU65PSrhzTdkzs1lSI/Z76SvqPMpHOhHk+E1PAMjq9YbxeDPwhWpKfy3PD1duA
KNZt0V4NcldFDJpnAcaxohVsfImYrE8+gEpT/oJvvAdpzf46VcHxXT5pedFQxL7Z
l1czuNi/FsYn9xXC/T1wy+VHyOMoCCnUg73K+zlWNF7WZDNjq09eNqD4x8rPRUJR
zk5rC6LSvTEA8E5RMZpFH2LhvFonahVUmz/7ZbynaNej9i2tqSELLrhjdUxAuEDI
wVAzr/Y9xcwdA0yZA0PknqOrnyjFCaSpFyUn0IhEpK90ncSt3z7c37eN2BuBQlzf
AScJP3gl/QIe8QQ7/saoWm7tGSFNEbfRpP3hqfD8ccjzlpSlB5CNIENbQX3DLHWx
+P31CKxM0PY7/7BubkoqdO6jVpnQl4MIQpVejxEayT39eO7JOTdY9odUJPyNPuVn
B8tKq08bwWItZqNNqsoeRh5KDTlzArtRjR9HjHuMRcjTR38npZ2sRHRB9r9xHQy9
gO165TCBfLmkYo+AJxL7RQ10UgDb3axK8Q/hL6YTUR69hYxTjcDXCl7L2g7ICwGj
2p/IwvaD6BWdwsRhcVJQ764bxYN1MbzJ8TaM8ERMCPWu5YkCZsIukkOow2TbUtp/
NuSpSayWaHOf/WDfrfdyOhoxZcacxm1Zq9GxWyqUyxtdc/jEnOZZy5Fc5IvoNFxr
qvIvpDkM/A8reCyOjwpA4UOR11nNCkzPgPgIXNgpjet5zuLr5vpIMj1b7n0tH60b
6OX/rwDWIJpM7aVCGT+Go6F67f6IeBY3gKigee0rjdOsnJT5TvDvDSJqgH2mUMni
d7BSjzjKctULm0YnzzBWCxniful+Krlf0ilTagdvNhfw4P84CUN0Z1Z3Y1abt0l8
lmVnOkrlDrGs4GOe2dOWxg789juxIVXTlV6mubqfinrAaEZytMsv2WSCvS1pze91
fFXjxMCkrggN15OKWYwoq2LSDmzi6iqgvV6RLn0wuzXViNyEy0hl78b7udzb74rq
CmdK+5eX1LiqRv+sr38dnaUTMlnWk2z7y+ajntCOU824Scd7XARE0IfYbFSZDzfj
3DrQUworydGtvUzibvwdh2PFqx5A9A/yB0W2mDQ08lElISq7swxQy8YdFKh/yC5c
IOwXPfmnRaQeyK6msZFbLKBRBu+3Z6EYshRLElLV6mLudpS+E7B9fUMgA6o6IR4n
iaMg8sxwMp6SFG+Hl6aQMnPeOQqSu1e7KbiOYvvDkxUgExlc/68xT1fRqPl8fX5T
deERYWHn93dFLf8AjQsuNh+/sXDPPpLkadGrM2M3MxC9gBzXrK4qaPhQ252BQ4y6
yEL7AcgJAe+BLqffIC0m12VkBBhJ96BijPlkHqcmCwDwKLz9R38nfpcve244wOK/
GTZDVXmjYZCqoEpWeN6ZKUQSFYVi5Cz7boYVYXex9IThtFY6Bke9Hx3u3YZxc0DQ
0l+527Krgu55N6ugyB0NBJJf+WatoLoezVvd+2iJnLf++SztxsLZfOOhb59JdCa7
QKaUDMd0Bzw6O+xeZI2MNNWOET+bU1Nx7qugbZlyTLlTLvvcEYZXL2q5kKKZ7qKH
ibLUt7uFhoXWKsptvRnWtVGNb+/Z2FxFj7mF39tWPyks8qdGdAKzyu5lERDMeJ5f
SMWD71U4JWtWZ+YQReGVUOpExMahq+NFZ4EihpVroRImIFic+ksbqBW5KAgz4v2E
Aj/NEQkPVZvRm/1qjlDoZ+CxXMb8OFjrrveIRWyf6p/swsz0kcBN24fZ8cbdCPCE
K4c15d5AeoX09QRn5Ey3ys05ERl6IU6gZey7WPO8J1twdrUl6YDYQ0hsiDLFRLSO
cHNCFLy/aG5QNWxViGLbG8QWMgQPpvaan4rCUB/5iAHcXXWyS9/T4G1EB22CvhHe
RnBLdhPabQ4ConPvgjKY649QEzUAWgEZDht1L5o8WXy24KwUHXIkLK6XOFiUaxHh
Xw60eYxp8WtyapdafTLgjOpEZdO5EVKlw3lTvNoYczPOKwt91RDu1xC0wv+Kuczn
ZheCHzZB8Xf4Vl8jL6QPGBCqjpfWPyl6422uZcOyBt8xQbkrxa9s44KZpX2AAnc/
o36jYu/zDrhQHnZjC8qrCyZZSjU5gmzRpQBnCZpf/d5urpAi6dOE9x5pGY7tWK5L
bR5bngmlY3xZxi2FfLbIG7jd79FP2+q6rt6oIctHTjckCjLOhO5KeGWNjMUacd5T
HXDMvPIezdsrasS/yM1+Kri4BAqB1f19Q8yrZdXk8pfgBXrNb6dkXCVWZlhIqOw5
Y3y5d6czRJqX7yWlv3z6mxA9gQvwi5JJduHffMyt4OVQig+K/XO4RLpxAbGP/T4s
g1ozjiZQ+nRrLJXyEW2KM//yyczvbteXH1LztWGNougWSzw0yIvu6bu0fCQxM3ED
XYMaXSEq/XF8nO0TAw48MUnbHJxzlWnXv/TyNU+7/O9DqA7i5Aabz9zB8S322xpk
bK7O6EOBgLTnF1fF7lM68d4JWwlG2OoSkNq2kaYcKR4gkD2thIPjG/KEkIAACARw
nUU0IH85BAzsV0hvHyar6lcQxDhyi+0swDAemakiH1fCxhooJhjYjNxu8j66yd3L
ckfZA59zMId423EKncIEd2tlLqIDX/4KOdpzQmFl5ais+ccg/z297lwh07k/vY2O
oaFWyUvkYIFld8/0fp+nne5vDWWeKPYZmAHq1by9ISgkv8d4vXsu1IzI5xIEfJeZ
oRZPqV0iq2YG78bytRYSMyn97IEZm/XlcOfgV0xnFxT+gErckQQBy5boeuR9iJUO
gqQnUJu88iTfunnG6mwcjmXRillK2RHJPlAa7Gxgct012/G/QccOwa8c+cIbIYRK
zHE2RPQiSbMOk60pSNcclJcNJNYHdAoA3kMiOjF+92hOWiXEYOAO1rquP8szHVzt
59+k5bKT4pKtysutySGteI145RXgoi6jmcYzXjb6ktiGwnraRK0dQOWfKH/7McLB
9K59GDpdyQJQun7bXUu8cqzsAxZBrwvtIYe+fRGxPIU54tdt7o9/bZeCXlIxZixl
0sZZjv+eQsLC+i5VjsJvOhs/IO62M7642UGtPLj3E0GP65FUkRgKDhlQbrfrQq8z
i7MmoD2GfC6k+McrnSZUEufQiweuN+sDG+QLg3+4pEtePSdkQ0W51ZjXe9Bx98J3
xFSrFBK3yGc7c4SMEYsN82dmKhOpa0XQZQ6tJM9HKlkipWH/6HuIPKSMsUF2Je8V
z4c//hnVsoOIWjF3o7zzXOowLQ1h8O+N23jm0AVyDfPhaijnVmVoL37vRIMxTPvu
VqP78vXzzhbPBkm36bCATVPlxDFnfs3MYDG3D8Qtx90ykxsIefaKhLzgsjPBBwTx
Xmh26EV8OZpQO1f903PY9Oa3qQfh1akVpdAwpWTSrt/q6pyYQQOJOXLYcljirJB6
xzsLdDrRZ8a1g8oXzUZnRztWsbTp8AdzzBiqGGgpGd4zHriUS1kMzeZbnEIMhHE9
YuUnWU+qOuiP5Gs+NyQxICZC1+zgFTY2vrJ1c/c8xGncmjOFZrySJ9mFTCocq8xD
YIqTTcaM8xZhSpKQwsaE+2UWQ0vmA6iK9hgGoAMq7DbPFmEghu2CK+O1JgqoEGbX
b2/TAwqLymRMY68s/jERkaJar+bN/JCmw5wcWxmTG8cDwUMmo+YE2nHnaq7Y3Ttq
6/RE74ncF1mb+t55OcHVgnJu5liI/f2o86RRnIyb3WtAD2Ve+jONIgddkU3sUJnd
klxwPB66VU8DzNm+kBJdXUPyIMprE9rfncCXyZwsLtxAz1kqj9CaETKyCY3SypYd
rO0cED1FvP/YjyMQ+cotyFzErEOY2RsoS3z3WIPj+HG2c0r4bc3QvRnHd0ZGzn/d
XDptDDuJgmklTH/LfwLGt/O3UwZtSYWbHH4vCUCSFwyLPzjIbGy1QeidI1NGV8wm
HHYgrThVUGsel8exERWbsEiv1kA5wQ6J78axa6ilKsuDU2BYuauOiBq2VenBTb9A
RrFIgN47R4MORxNVSe2LYjRBVSgH9UETkyR2yk3LqXmM0FS3xbLZcobioKkpmZ77
aOMmKf11HM5LkYOZQQiUD05gtEX8Zz3EkZx/QGxP10A/7e/+NohXPSOGoLPb2a1X
fopJxk6HGqbFvTDjirO406wFpNewHEVvTrrVN8Kv9Ix7ZTH54FLgGhY5vgE2IUM0
JQH17SoGjMFYKxxV92z1K/R8MQOXkFGfTgSy5f1MvLFS+m6QzGwhzPqbS9evwL6N
tY9I/qLi3MIf0LTTdUkWxFoQlD0B8YPi6LZkdxvT2UHndBGBCGXfQDgGBmqoF/wf
nqXojWDnHYUAn98xA8q4Ran2Gv1+g/3U7IfadjGqAXxGqU+hjk6RTcLyzl3seXqz
DbdVYYPKDD7CmOp5IyXUGnIYt5j/HcQwCD6ox1n1Zkw/xpR+46sZE8acAPHPqFYc
kBhcSFqd+sJlN6yoxlL0q0FDov6wXRjgmyXDHN/qhV/I6qj9DuCN87ug5BsJm40Y
jzKlRMPSEfmUs0jj7qvOnSxTj8hQwkZ6OXcE4Ls8uWHx4chXI7ku06SyYBTGrNWk
+mDjBSd9LGSSkFRnV4PQxG+N9tIzUIFmaJZGhIZb/WggCCUBe3lTt+2NOPrnBWq7
fn7qpzDdF6VQckrRWRkoVOAnpEbrLTqcF1nbURYP0aC9wgYZVM9d5Pk1JV8U8dLc
9ds687axOTcvjm7n24uAK3K9WE8oDtFanfcuTYG6jILrYAaoNl4nrDRDkXVI7W/B
KogUchBFb2W4puOsjZPtWYPNtQ/8eQij5ZsBOd/Ct3VWOh4sMIckKCInF+7MYwbQ
xwk4bJP7U0xARFgtX2B/yU8qX0N5yVUGkNMvmz5eIRiWAcrskjOyR29wjxPaIX8c
+uvUFHBmQj75k3/aQhhsr7tFAY9HHcdVTayyXifh+JulGwf590Te91zdSjP0XamN
deJQP3MbXEpUIElc+OML6bpNE912my/J8Z9EBr07vvaiz2jes0Sfvw4A4AnzAkmh
PCgQqbyc9PF36T1jkXmardgfnRp/fVDsmnDtkwWccJ13D1QiemYQLwb8aq6FP8Gr
4Aq5N/AFkDCz6Iq11yTlMy/PFOr8WZiM+3wmCQ2gziMy7PTAQaO0g2bW7ZgnRvSZ
UIpiE7nlK7IZivEmPqUZhavALa3Lv0vnIDp7gA/Guse4LmlpzCNohxj7WvjDUVuE
xFtnlNf+oiQVnWQai0JdLXYJIPZ2ojmiFVXppFeKy7PM+EdpEeO3QN3OMxQf+yPI
hrgtyA7s8pjmuNyz/Y45QKNTOpkm9Cdw9SpA/FZUxA3id0TjMBhU5cbgcNkObeZx
UUGB7QwONz0VLnQSStyqdPDpLJ5jEHvCDi5hoaITG6IMY99//pj8ecWqnIvDjDvo
tcVmuyXjB6dAzXSCX/oEzb6gelkWzQicMRe9beEJwILFA1K8lvX68eYMo019+Ojs
eugleeK5eEGS637Ms9T3K0gUdQcbiyMgx2LK8G9WfWD0HyfmewoZ7Q3Tx0OXrjGA
7GrvgoD0wfKft6MMA9ph8X0RetEeU82XX3q3mACSQJl7PjaOCx45PATbYlUWU2Fd
/H+B5vMQ1rK9Ogtqjkj27F3oSSkz2O7KS/P00Tg1YcgR+RyzcuQUyNKsKqgBkNK7
GN45dhuF9dFjjvhUfjnau0lrzUaGvJr4vM5A7xL7v0eKXZvPFhlYbpdaa3ueIuZG
ByUtWHsdaWDH6636el9pOHq7S2XslKnZ2MCaCV7uslh2raE0/vhMiUNbApK6/xi6
mNcEBEGSzefFDu26JycwaPLMhe1y5qD5r+0VSPxTcyjzk81Nm/98MWafp9ALXdWX
5V/eIb9pWWnAwHvG5WrYvI2HjpE760EjGXBZmJK6QPO3F7d98HwGvGamNwuUfPDD
4zEIJuZt78H2r+lON3VsQaKcy9n51pm6yPP7UB6s7C3ihwGjhjfWQhY9NIju5Oqa
gvNR1O/hn9i8uEG0/g2dR7ymhDb6WV6fFQr2uVDd4bXTSDvJuD/lBJ1SwEpPuXUL
toilGRpUBz0u8XjazUJG/5EUQcTIu/8/DH4g8+oDl1E98s3lwdMG1fkKoT/dw2+z
yBpL0Q2hUWFJkr5EYXCDmg/t/MXSXkW+qQhWMXbu2vXcyLOlOcxC0bdqnHPSYurH
7PB9Vgqo6CFEG4BlaJOeCQIZlPdb0NdNeEIeP/fYYoDBWRQgPjw25dUnGwPTdsAm
LZZbPgdfgGcfE0nzXjSSrUia3gMbJ93cHfnVL+J2uEIIXNw/kVahiT5AZhlD4DV7
0q2yQ2MO1vqSOssXiJtrQWLgeuhs1NiKi90CZpYy2T1XlU5c8HbAZNMHRjcEpqDa
y1kbHnYL5pRhT0erYrnWMJO6+3C0Q2GMKT/Mo2zm3T+OGgz4VV/Zodd40NJDkBmF
yXs1uO1DMsLD4qF/tvXTk1aXHz1yE/CH1zO/HOITC/USNLbVCif5fHMNym+kCG29
20jOOljKdk5AauiKdWLxbMFIlfbV5f6Y+uTScmHjPuXM8xBpI/w6XbIlMXMA39HA
njBCzwMG17B3odMPlJyZ3ANbOswigU6YB059gvuF+xLeyCdnuY/9PEGU49jpAf2Y
iSbBbU7HljzM7baj6Dv/s89vsgwDZrZTzzgdSxw6XA2dNdvI9V7d87f1a0xs7dEY
/Qvw8BInx8LRUrswLcQHl4qvfmMQb0qUvDKbwm5DLQbXwuD7os0jTuxR8ch9lfA4
tklcaSC4AjS7v9IneNt+4269QovcB8mRlISM/2XPDjIY/lo5vF41IrEBAo4hqI+F
p7zR9EE8bxtBADHX036sunXhPVs313/b/YUBfL/L07btOqLbSW4APszzsSUMR+Sv
i1rVlDPSQ/msTK8ITow1W8FqNXEfMQaSqJgRIXfEy7CAgD8N3Y0JRDI6pWAzVyqm
vBzBPqGQeuKFW4LidrLH8PbX+pbaY0A683/mqLD4KDgHepAnz+BWsleNXY9I5iZ1
q13il88T4MN0/fr3f+mz3K8zWk+MdoUTiXsImPOsp8p1ItjH/C1lfss6qhHuHqLx
xDVDDWq/CiQIsFi4BqS1MQfMghD+++D0zWoMf41VwQmA0KbOy43tDt76Ufxdgj/8
J/IrnFi7WQWqc0bccFQ8agoe90zKXH97i52cRuM6vQtWCUW2f8hSHY45M4YDmqiU
i8y2Dp1DW5LxwtnCuesD5Qpt1dJtWxo6woKX7P3O5nxsPNXBLkTtNYd3ITVa9ikx
d2M1ppxRXi0JdShIAUfXijS+lcoY55zyPcronTMk1n2S+oPuaAx8BmfKCLp14Zbz
rTm6p1bjZVagCCl+4MnC6fqlp9PBdPV+sVLviV7tkWmF5IQNbBaUAooAnfkvyxsr
tKc+awvn0gm8htqdQE96MoUzXyvCWtWQ5kN4WSPgOy9zbic3uap0KhwkmzfWWPMS
efXP0NK/58+SXBWQbRoB89lZlIwgFrFAV/q23qrKV6OGyO0a/qWQIBRKxA2+X+rv
cttrTQE09o3I4mDj8CtVbjH0sXmZ5cQiR0d3O5kSqXlqyT7yCFYb88QAqJqKpYu0
apl0nlJzJU/4k8Ld5e7TKd51dX4vr5bPdMNdg/uvBjfMDN1FLBCd3s2mQLBanIin
07M0Dkgbv3dnUaKa0sh3IKr0PD8VmNJmlm/v0BZ1fIBrw4wRBLz/hUPNrhULkHH8
CXrq86ADoT/Rfd8nTSP99+V8SBKbsmktnGlM82N5W6DaoEpsQewLouFsECgVu3ms
VBh+GC8Jske/uAglFeLeuh/ksUi8L1tOxJS205nfgqH1a3UeVJEYJXl/dPRa6lUl
EXBfQXYMceyWTgXKdl6huDL2pmBPZkqD2HkBTsRNOOKtEeKXDDAOn7sITpHRtxRT
XMIfjZK85qwZ2eNVGuC4rhyj36GQsBbYt4i6nU3KLdK+XrLcx6O1LPZ0yhM+NTlv
295WerQ/8DmK4nh24RoO+/Fc5F2q7jXvr142QqzmvH2BM/HJSyheN59G07Eonqiq
eTE6a2H9ktHLuE7VdqTgIiU+uCDd4HgzNjIv+BMe2qm5NNdSzSCE3yX/wBF+hNeZ
ycjWoORy+Kp/80kx34Yn6BrQd7LKcYEG2Rg5+rfkKEOpi+09i/wq/aORBTgJPgfl
OEB9gzxs1VTRv6c1bzkIfyOo5mOd83+NEK8XVQdUFbBKZ9dV/R1J0zYIYFcX2Omi
xUQJy0hB0/VEwR0vl9K2xTC7SBX5nnq0b5X7f+HVqezKRhwqcJ3Usu5miKlNeCAL
Eeibcd14yvoCRchNmI85HVcHgzr5PH1hs6e3JPxqNBjTrrJKdvJSAosXADvfyfxn
RoYapqEchfTPDk52mWDbG/Lck0r2Oplr3KeIJfog8Ck7OBbD1G63ZX0vU+gH3dec
Hpup0PkDc9gHYN6JaT3bRqQBJK1QtHRC2GjJSCUDO/7KpI9k8zuzHu+fng0kDXWq
n8kwreTSOJIMI6HU7xqqGZUNzYai0dAue8PiFMd6aTsmLUL9mz5cNoTq9kLhs9RJ
TuC5gJwPtnr1NvApcDmexnpNZvTCK1rOIW/dPVFLpDF8SzARL9Ggz/JK0T+fLZyJ
slK+XZRdXafThGSUevv7Mq5u+an74UIye3SvTw7M5kElWU6V63wLI5mZejeo7qtY
FZEkQG2zyQm0Si+qYP0zYNCfMIAqG1sbEzygOU1o+cYIGKdjnBPbK2IbvCNoQ/v4
OxJ26FQVxqP4gwH3IlF9m+9H2pHMQsppa3liGHvyz442InjS7x/ndO/C7CJBvehP
tIWiLRzxMf2KIlluEzUz4j8ZkPKuksjCrjh9s+XXy+xEMuVeAM9dtV0mxSiqJZrR
6XBm7qzfHKnh0LJYCCkmQ+AHR1hWTlnrVHM+5YiqfzlQOfCs7A8jSOxS2f8a5Kpd
IYtx4bGYtgyHoZC3ksK2vnLo7P74coq5hY3xJLuJjiptY9JQ7S89SRKePwYrkBkj
tVdocAm9MHWe2Q875K0hNo+7f51KHNRL6ZAF32huOHV28FrYarMYpZCwHAGtjqrE
vADT9oZMggqMxECQNfigAS/lZa7ElhHb9L0+hggJjHOtKnCd6q/qGx6RUZ+tOvH2
U+cRB14nOjHeNq41aD3UDcLJVRCvKBTjqNi0cyvB+OVyO/ZvYKJ+c31kz1bHrrFF
fQeEJLIeWva1UYANvCFm9/h6kSgLfmbduZAOYL5UnF8/8rmqt55ltqOrCLpvi8IG
GXRcZ5/uqpylAavvezDZpR8prcL2A3Dg5i73zjKU0bcWAhSqnXG7Q/KII0mRONyw
TH3pwn5Q/7n1oNtgg3SMaXq8jUFum2dOVtIyz+S+aXNpr4EJwQaDkzWL88m3s7Ur
Z1Vb4nMjir8J4clSUCd5p1MF8htacuAkT+71OzZXv85gaySVGAwOeMvvxDSKuiVJ
JkPBESoUhQp6Z/sSZMDh5iaOKrjyepBr2djc4HF2SNQPUv4wocDn5WOwtGBptX7d
liQRwTi9c+12jSG+cFwRH+SvVgDlGtRMZfj6AzxhkaE90L7D9xbAZjzFqOlAKgIj
+63KaXSScOdIX31JAqRUx2EvR92uSz0lo5em+/vmEib0N0rezqlPBsqebbcmhnGr
wgROadN4Ep2rJsRlEIKp/GppatmeVFUScPnYqkGetvWAlr8Z4/zBqHv91accboTD
t0IMTvdHuVGDxqS6s2RebBbCMSrITGcQTtudSBQ90+VRMFFWe2XbK5V/H/0tfQG7
oMdfqz9mLFjpW3Hc5rStjgrOw93omkG9nFvRU0PbgDOhnn+ckl654I7M3YUw7eZC
sM3xQIVMMqU+G3e3/MycwgkpPdgyNRUT+167367UOOXDuhX9bsB/v2a1SNfFUG4X
gnGREqmF177YCuYImVf1vL0k1Xvju/ppa41hknklCpkCvMmifhD+d78ZMztqKkiF
PMXNBvxotbYdrg0BD4cD0knj33LuGQTbPBpXk4a5UH8T8e6VIuoT5i/DLrj63t1p
POmay8MP0V9oIG88+2oUlplhekSZlZtWJJPLCvt38hxIKiiYpzSffkrJTo5VtdAs
aWAq7zSbRjp2MSm7GefYySccMWDah4mVUvVgGZWZqXfxEw92CBZivvROAau+H8GU
OKqZlRmtO7V7RzEl68A65EKor8BrTs+U4KSJgULW0SFchuKl7oaeovIQsqyaW9Aa
gzdvaP6V5GlUQMqXfEmGaa/ZXXxLIFeDGVMUCsltgXBstvgs0nk1TaLo0CMYuGh9
+G9wkG2HpeYvM9h7RbEywcxVxn3Wfopxrf7XVtrc0itzksIhTq4UMflkuaOuHxLn
Gsyjl7Dnq4RyHZQnvx0I+OZC/8e3wpXqRPqqEOM37J1Fhs0QMZEt1tK6vaS619s6
HXGtnp94epei1ThaHKmPkH/RndoUxJDoB6yQsFplcRMd77C8XfvR8pkCUKxSACZ+
3TCpAg8JCUmvtkQnO3imVRwTgv6pfLHGob5vxw+ocDi0v/mAOosIE4DLNVtBmlx6
mqy4hg/gdcF+QkHf2G0OVMzfZ80zBfb/KZ0lrD0JEFpp3733oG6f3MZQtn7rGGGQ
TtKMBdsx6qxFqBptrkgaM3soLrJJfwbYivFm2cxt9kuqafC/thMm0A4oecTUceoU
mZMI8KaNaUXq6MePxheexeWb8tzTXaHA1F7O7xKjFr63p9c801K58RQ5L/Gjk4Yt
/oBwqkWOd347a4JMYnN6mSbxSu+trl543mwf+QUoJOvxb+cr/iHTcalCJ/foJEp7
eBTQ4V+nDTyHBkVh+b6+/lMxhE51sHR1gwqZkCIZlzxJkcyQLGMensVtuJGGW5Pb
ByRQuWiPXu3H4V1HVZN0g9mvbHns3ZUdwUeaTap4hpjy67UkfyIcMCkSGLHCyAXw
YwNrpzJRufWvp/ck4yR6V9zQkunRjG0GU4iInZ7ifjyl/aYCHzLpUgYpGCT0XtLQ
e0qVW/a4HZTTYx+i106YBKEiN01pVoTAz5fw475EyIvD3LaFhWTWmiXekUAiqCuV
/l+se1zALH07GSYSMTjiPnK5rFg0yw+UagJHWC5rqtp5kWrvVhL3e0EV8bYNIaY2
/e82UYtFjzj0YqzsPePswarPgTbfsRdJUsRzTSp2LSc32HKRhzGVsYKsaU0E9IaW
piEMVbg19DtMzr/Z4XeDzPCeyavFBjLTb4XnFwqJTiCQI/C8aef0LfupPyBrvNoz
A60SJJ+AlgqUO4z8xhpwCNNDaU5audMMb07R3yBxMUCTJf4TmldJhS4Kj3GP6HWs
rLwhaTyc2RkdYvI7RrEl282Z2n3ngdK+2IxJoLz83BqTStyS4Hd6lwTj6Z2ksHq3
HYsSiYddk2cPNSO2yaIxIl41J9fXj9oDN1zxEfIqIoHnzaJ+1krPVwB98sxIWnyh
kjm4TrHakma+NZIVjOyWaZPBCkxRO/m2T7SWzOe+bZbrxXkjO4/Fq5Ilh6H3I1+v
4Cgf0iEeQAMB2GNO1YN6GtILTj97WpRJSJdJas7IPXdVW90/9AK922SdHaJOYTju
FziWM2xUMG+YwtekxFctHviQNt5vuMnDr1+1eIAJ1STvGFHUiz8pQiMRmT3QoADL
ZXG52fu3XFBg9iMFYmJsqnehXUpEHXQi+uGkqrY2Hfrlz3VXf9b2MmDs+woGNnRR
C9yiE7N03UkqgYVVxQC8KUKkE5bHW4Qj1/jUKYCbsMyFex8PliujhLXkGaSTqO5R
xGxcgMUkDWDipnobq6uLEwbsLnNiuA1E28zDKiYnk00qc539gApTr0eQamY2J5XM
JEDbkZefoFnV5Ra5LHwWrYRCoVXIW41YsLKUNA0WQfH9vWLW2KwrjvZ2q0Up+5bB
mfuup2LbtzMn7Rsr5b6Hu/3rZHW1C0CmCZdyWG2UwUWLR+k/LEOoLtslhnhT7ko7
R3hmwCxaYRf1Z/QDbb0C5szP53/qcQfH+hIMQSRTW1PNw7nBltPLJFgVTfFDA/D4
U/tIGFa+g6hnDku1e5NtIqXIOtTtU3jjOS/P6tSExzvzNbiTM5gK+A1uHcVFAq8F
aNVopFKZMpBB4FECDAGzyVUZYx4zq64FmfjV1HLZ04G6fKr4ozF0CaImO9Yg1+S5
Ngnwag9yLGbe1HrBa/qsA+H6Ogu1U898gmpwFHkWhk6iXfHjZQSLW3K8DOXS8d5c
vQeVugteU+f6Ss/vMSG9qRFk9QgSpawNEGvPAipBP28lkQG4kYCO/rQHxyEEVMte
E3laF2CWxfxZL55gExQqVmrri9qMY3LAdiSI8+p8hGL7bR32vQ0l2bfh5y/6foHd
1YYM95xQ9ruVVqoP7qFB+YUt9W5tYKhmMD8TByp7GSchL4JjEK2BZr0U/L+ZI6XV
AZwRtr1mrdoOlfXcr22g3wuwoVOwotIEV6GlPOYee2Xv9llT8T9QhlAg2dzJROVO
FheIdbkNj2mjgtRCl6DN7fJ6NqkoWpyB1KBXgp6sU6aayEDuN0e0XkB5LMXqssXT
TD4bAe4FTBHcI1GvYjUvhq8UMSbRrOX9sN0TDdJfUHxm9pXG6PyU/++614bw6iAd
TNbuw8lSozSrljdYrZfdQO1Ax/B/1E/ZjUdwwC0UA3q3JVCJ0V4BeDgKzNpPUOJY
NRzkEFK7r/sLsi5pfBhI5H7sDXKK0PdDluO2gkDqxnhqNeeXpdhLAaBi8mgkhraE
zIJ8Il764Lz4CCZhd8DteKClb6IZjIU02f5BuQggNe0uIYz4d2OWTjlxwpenz4Ee
EM1OmeDq544M33yxb2VrYBc5prOXzBZjaVkpwcuCTW1bEVGzlkgJx46t4I8PIC5B
vRidde+tNxu018Bj7agt3+waBOj0VMQ+4xAhnXaKokFWtOJ7AFHioNOQNzfYOHaY
YfEphriqhHHtwepTpUTOXDmZXNx6JrFSyiSLx2SWdiM2mcsx/RSwLKCdpgpDw8kZ
pCgfSQtazFaLvT3BKHMgAcK5zilaelkNfGoMd6o5Hscl2PLBNJU0B5NgKlGSQPhW
L42JNXa+Vz72KHIzq8om3U6V/1AhL/xXD/ARyeMNY6LctaPQz+MkoVb1UiEPP8U5
XmH7nTJBVNFsPo9rb6N87tGkkIgmeXtYyGHkj0NMO+BSLxU0KyCNTb1NfWBn3Cei
UVto+ssCLVf4jEq75bAVYC8qkRu/sBi04JfRhIV7jskFc46S6DKoq/IAmkvK9lHU
mNeloTZcB4i34AmOcsawbQW9V4OzN5C0E8pjpTvVr011YdRdprhTHb38zXNyL0yQ
7+0mzBAqYNLhIKnEVgiq/iOzPhnDBVJrx0MtavkUaM0nbnqwdOPKGFbgSVVoPRqL
t7UoMjXunr++SCTZ5wljMWljtrEzKKbWZmTaeIYlx5+ID9f5oiCj9ZsYCbwr2W36
niL8oRK4LLN6+4QaV3b//BrzfdqcD3T4RG5hioZRWjcFf/BDjqSFO6xe/13VdrZe
5VONZpkofyfaFAxaIP06LNHLiIvh4BQC5jrV+h2tZDBQYdJAOeMMcMWNeQgGwbh8
Gi14c3Bu/JOYoCntGr5491E7nK+ap7MmGafD9TYlNQ4B1vwVv8kAVTPZV5BjgYZY
syv3zjzWwzdpq64LO97iPz2FPfGy86E4wlhU+kHKI67/H/HUeUMJ+hh3CbvURcDb
BymSSrMBxBVE0hM2hnStZkaD18CMaUctSJO48cp3ySX4wnZcV6PlMN/6rVZl/kBl
fsFuEeF7o8Qu/Q3ZpmHFxhL6eIk2lW7ozIieOGTLopDGlatMS/z7vGlM3h+wmmh9
9f0/TEiHb9KSEj4CjCANIbjo3E3zlS4oEgh/znGyT5InL0Ec8yWRgMy8emy9hQmj
7h3oPLj2/9+loVl2B+DI+S+HLUpdGZjYlpxuvSnxooZEEGzEYb73iVZNZH6i5s6I
VaHHkCJ5ju2xD0iGwR8Pinf8RIzJBic0kDARGc99n7b1tsM3nHKDRjawrNUvhlZl
xvLHc2i3Kv+tFxYJa/Z22iKd1zaRInETdz4/9ZZuCgUnXpImghJdeL/Q0fE0iUXr
G1JfpTQUfDEsYHObb1vDllYeYcj9WCPxESj95NLti+8XEBkPasYBH07TzFCR8jb/
fIivIJahKcPcnObgTFwRl3sUCtUVVDf8v4v3CbnJO5Hg2cQdJA8H7En/6Kkyqudl
76YiA/HwOL7aSjElU9zvhRKqetdvYcLqt1JhFVyHkj7Ck3tuEZptlRpFNO2YkqB2
bk+CmBaqb5jkCoDwB+n5tOwTWCWpURaatvVxqth0Nfyo/LUfUN/Wwt2B8hcK7HC1
oSGA7fnihOE3KuAltwf/o+WEfW8wxMHTA0883oGHZLZHp3aQSHIQNLofolYXpFv7
NlODLKE8HTE0ySkE85i+bhgURFyNpCcSzDGad5S+W3CGI374q508L4vQhfXyGhAX
Rv4lv8X/nsTNYXwHcuGUVw43Zqy2ZSvawxMk5Ek8r9udUxZwZctGXU5SC+zShM2x
+Y++mfgsW0irHJvYMFaUQp08NcfDVVos0tabYrK4aAQO5CUkqb6pPs/8DW2WK1tO
Ysd7/t/gO83W+eMyEt0onqvwrFh1/Vh8vscm/qJmjYZultSppZqhouBb/MNtgLvk
2MNredyiiX83ewqxwz1HOAGPzDsHUe2zZ9vmM4bgAAqaSlrSkxL/BoXapINnfak5
QMmWbOPHiHPuDzp/blV/aENwD5qBgsiFX9q7EMRRmpGA0v3em8LEFyqVfFhLhCk7
5liIZymO48n2Y1anDK9jt/kEzwQ9xGaAjb8ErgbGKuh+7j6COagj+tjux0oE8I9u
5Cim9TdPI3XqvYchUbk16JC9jiWqh1/uBPFUpWTPTxxzokVh42IoDm4UszO5hROu
kukqbV0C1Q4kOX75sF4nWP1QJ1YB+h4tw4uXtfutU6rOoJXh9uZevwSEKh4huyPc
IlPltdaQ8TovPrLwYmleyP9q5elu6ZkwNjrTCx5knjN5sKQHAOlCLSVCch81YnY/
ZqMXslwcBy3QFl6RQ4Ym7LSibK5cCeqQQtcdTzhPG20Sr2CuGOz1jtls9uFeZzbP
cAWkgVSN5b44/+G5l6TEQL9a7z9PY0Oe3B8tuHL9e69r4teDMA6ZTZEx4cjuk1JE
xzdyK+HAOGkSCAYDyn7WeMPXYEKh8KdLOCzcxxhx7Fc+juiGw54nQXRcjCsijyQE
r8tIrST2FDWynk4/nxf80uzUuexHmTWvjQ7KZkocfDwWGphOjwh/rJT9jUtD96NB
3Sxz9xhjHZe6on33LLGR1BFLDDfWyuovGelV14UzJlCcYFKPCKi9I9f/e7Ju7b1u
VyZmtK4FLcB/OaYO2LItjVeywbWfRzUIANQxvekcFJoIn7pyvNqp1MTYk9+71xGh
fJq7A9kVqoELQaf5XYDtpTzJmYpdaZX+of2Ud0C6WukiH4lok/7IHAEkncSGGIp2
qb+qhsasJoChiMaXTpSOrwV0Ci0IrQp2Rixksha4P7diGRlQQcK2hAIbXxU/3Eoa
G/0UZYgWmv4Glh8Lk4yJrwy5WyY4VlubqEmqQvo2anN4AGm495+V76NhOOnM/AAd
81fx80GVDVFV4ylRdHDgkWqAx8OVIaFhtxP3nQZgiBHAny1Hx+LyQXZkGUEg+TKX
ShNgbWU0Z4pciKW3zA329j3ESm2sMvl0Hn0RVR4qlvwLDClZ0VuFLpxwhm928aM6
J0oXo/Xdj7zVf4KZaBDyPY246RfDGSoMzLvNF3LrpFvEzw9dmxIHaUrf6/sjdxWm
Mdc453CnvPO3RSVAxw2aqHiXrt3xRAl1jSQRHiWcwpIO05+b6XX8qixini7HfAZR
1vMu8bxiSsrrURDsl4sUAhZ6moAAYDRqE1JqXT87xmVlj1SRhoz6Z4VT09WfjUHw
XbRxcNGHH775Y5LCye9VPcwEfWP9yuwFL9vL0LS9wLEq4xgv5VDyxSE1UsITCOIM
8xHiusVIB04gUxrP9ru8Rkx5Srbp8HTsdhWCJ3kWx7V+lOmd5LLktyjkCaY6OQYe
S1P5RLAX7euy9BBjshNsUQ580RW8anmy0miSyKuf0qiAFvkJHDNjy3g2QSdWGM6J
oLvY7GKT6kEMaa/iGTI+yJaphxZdgt7Z04XN2fjkTbiNL1PSC6G5O2/i3PXgxWeo
UvazN7qEJLzl2zP/FxE9QlYo9SI+NFYYQXh/M8VPghclUUHo9gqlodW26ScyMQxF
pNfdIo6YzY7SmyCZzQKP6rUdIqX/995i9+VA8hIMU/rj571YEumdqFjHV3zKCDcZ
Cmpz13Ote8JuAxJwPvGlShVk4mccdvS4rI+fsixl9bPddm3NHr1LkR2/erOgYxJ/
EJwMFb95nA8I01PHiddANhLpx/91x6lH/8G2I9hdMwRUb6dMoYKouxiMaJ+YgB7F
5Kaem26uU5/EV5bNaP1Kw+2etXGCU6M4BSp7ETWtkT1saGuugchJevn9Jhl6Qm/2
BHoPnuFZeBufobK2NYTlQc7hb4sE13xq39oT3ww7whxz+p71y5wBQ43SZn+pazh3
kfGTOAeST8OKYJZIUi0ouSfqEjypuWjvF8q/dQ6h5KuYWqsSJt/kPMU0NgYVXm0O
GbZX4g7Bx83wa0UkBI0z41gvu4oVOzdou6Omx09TrQgt4xSEZOdHWcDK7XPp7SI8
bRRnAgMt4dSHHH2UJaxxhT1CqExGs18IsJ0dD7MR3MP/rFafc3QRFSI5nCWnIq7G
4bhbEWxHshjjtPYCI2RIfUtGdFpnMEAYVQ9RnglKuJgGNyKb6zhevGCfLE78lty1
Cjdir/DK1Y0u6MXI8spBvEpPAWs0Yv5Y4IdUrX/TeCw9Y6m+ItabFrWjdvXUBOU6
aloUia0cZaOijMyVSa9r+7YIqSFFTjb6BSobIKJU6oyG8T0wnVEJS8pjqV01IrLO
Ped9ZCWRBaZKXWenVTXzAEGOmt4xXOfWpw+xdXCyhs4sIx+PINm9sij7LyplwCND
rrg2GZNcGYzfp29x9rcNAuPAJniHquMwnMx1USgTbQjlZmpyOMO93WMYbMTLfZj5
nDljZPgShnn2grzWodNoAblaPoF9e6EOcXSxsOch7iksYHQ5pDHjtTTKHfISIFii
PQo1Rn+MqlmBEwwznEFn0WtQKwYL/arjyzj2Otp1lYUZN0+092/PaJNJKuGdNDVD
4U/uWao5945CqUuNZ/8aDrN6yoRdZmMC+0jf0fj0DCZisAC7T8vSHRx0yIKAw6zb
eYGmItt+wMnq2YbmtYIjnEjZEQn3pUJ1XBLhmcnZqp+TBlPly9okYjH8uTavQdbx
vHG5un4xvADbP1IDJXqbDfwnWt0dWqKgYNvrrOWtSzl8QYNvHytLHhkmUBx2/Hoo
RWmFIdPBmWT7xfTbSa73hU7t7Vx2eUJy1URrsa5UZszsdsrl7hMO3HlfotlsWQv0
Tqv1evJIEXa0dMTf5jKkaACJoT0Ho7LzzOtyJa8YLOt1RwE7ODHMPzvBiKkHjWIO
2luaxBixe1yVTAdRws6xUDsEvGAYOgOebvBjeSAFTHzeVqxdqmZVn5fwTWqMAuqz
mbz52OFaw/AqwiyDPxJhFnj/ms81eTRp4tyWjnHMhtYqT7LS89gS0dBHpefWEZ/e
pwhj2A4O5NRGwcBK8+HI/IbtRv9Rw3U2ChU8Re4I87Ycb8LxNi5QuMccZUQJzx10
nY42jctMal/A/f2fqO6hS1XX27HMbxEXUAdPlNUriwVa7nyDerbodtB4WcoHpJjn
g0lYAE1Al9etVW1IdftgclEc35YOV+l5RNrFafYUh5LHdZQyUB/ukujw2h26EjKR
/sKPpbH474qIkDhh7efNd26BIend39VYQoMIR1VZdM/4ItlMQd3LODAgzbKn/Uv7
bVRqf9AcyBgQ/K7Vr0gOuWgWfIGo4l+mDPapyHefhHLy4DmSUZ2WwFm+6Xpm17VV
yYHK0pHw8z2oO87qz5vZLZuQ4jW5RmCl7enMG7OCRWQGJpeoB1RZ2UFo8ms/XmNN
B8QiTw+y71l5yuASuzv8GPBYaelMBVuTIhMPe52f1E6TPqyjDTtHle1hJh54gI8F
Zs1OmPhXMTWwg5GprhrV572p/0E7KGm9U9eV02qfYBYFB+4Z4qIpKBUXwom7g5fP
G0CnSw6HLYqI87wY4ax1UrYoM1GtIh2PWPQGPXPn/OgcNue7IU7gzi6AVudsbQ6U
+zvtRC2kKOyyQYrXfwbhlNQlltYXSI/jeOUz/6drcdPZTLc8mycgUIOhXAQkvrRw
skiOH0/nlz/LaD7C3FAvcA==
//pragma protect end_data_block
//pragma protect digest_block
M+fCgWdAbK6xkPtMoO3IEtoYT1o=
//pragma protect end_digest_block
//pragma protect end_protected
