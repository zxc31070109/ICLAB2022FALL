//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Esgy5jVOEM4wr+ikL9WubcirqvSldnsPzJGV5Odxdt+rqCtr5AG8QDASVwGA0kNm
/61rn2e2m6dARBI2YkB29cq15D9CAR7OGh10o+G8k1WiLVOvM0XGdt1mhkCBK0bW
KnaFEBD4qqoIvjF4wmANPUWDH8cvX5B/aha+DGcTkl9E9PACRMd+NaKnLYQ9w8Xt
iz+HwHPGr0sgbmoHZbd4UDkrabxA5nRSbNxecRjjIHMjrnL+V+RYkxlODjXi2Lcy
7XOfScGbQ+1XksithOJQsj2vpxSJt0fWmaqHS2Gjt7HDRyipxl3ibXNI+WzfW3UN
tKiaX0/caWewkS69yyCvTA==
//pragma protect end_key_block
//pragma protect digest_block
DEGnyLnyAF8QHuCQF+6I4S4X+h4=
//pragma protect end_digest_block
//pragma protect data_block
5i2UPbyK0/mlfjJpCcEbjY2wCiQHfFMpPxhjTKPBPH1Rb3G/6rtl40nwpz/DCTEH
ZudEm7B/zfI3lcJ1CSF+ZCYettdccNERvF8PgicKdystNPUbRYZPDR97th2aK+CQ
EfM/HH3tNfPrF4kIbT5+8HhPs6qpg4NwslS85HfkrBeEGef4nsQE5gt3rEZNWwyz
Qc7iDabhq6UfAgDwderaKlOOgCvHiT0EFpmC2nvakuZxAhHSl1vjKJrP2uUEs2tp
p9jqfI//1SzTXhTDXnZPzq94sealCWWSRQ4QyjPBpeiBWnaG9AHayAwGdZAzJ90A
vBybGB8lAJj6CMrWAwngCg==
//pragma protect end_data_block
//pragma protect digest_block
1YVAh+n/P4hxVUmKHE0zkKxFJkE=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_FD.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
CJ30kgi6XhUMv1hclScWAXsrsYAtUh9GLmNKdTeklmYRuRZkySSbstsuC4oT38xc
6/3r10V8jTzN8oqF3JGKZEIB/U7qOaP5p6OrxZYTCCjm/IkMoYn1q7QGoSOu9+Hp
BtBYEp6CPc//xEG8P6laJlo+6+zFkWgGe+U08suUK+3Xj8CHxFHamjtpfelEp1Cx
WUgoXGg+2/CQYYnvLm5mFaPpdPwhQDV2vP2X3zN5WDxo/uh+LRzK5n2vmrJSwVy4
mFYix2sKPpqjzKcdhlz2C7r+WTDH4gmekJDG9sEyUvlyQrO5gngfmg6RBDCLSHhL
ngze2qImtdOgR/WXH9jjiQ==
//pragma protect end_key_block
//pragma protect digest_block
L62ATVdMoPgLhSIVnIHycfKfsqE=
//pragma protect end_digest_block
//pragma protect data_block
5Y5gFAolq+sdeG4h3lZbonkWpPDKttSWf1tcRikpCPd3SI4KcQbapeuXooDemgrN
JXGb94X9jybOdaifQGAhmmOciGZ90VVCACP5GT3jWtOIftCUSRwuepFCUxRySfv3
I6ptMcv/wP6bq5pC2/EMeVzQ/tttGUH9pB4cR+S9nMGa1+X+VN/OBejzyuMyqOxg
F2Uf6lE2Vt2XWBe3bkWnSN3rq6RWrLZEetHLAhSaNmdZTV8MYlrPEA9NqrkmD6lw
l80pRWZWELalIxdbROT+0c0SGbd9vgVKyyMUHXX0IIIC3fsozyK7VW3X+ldhrYhY
2hPpNPQRSBpIGM9nrbqspTfaRbulxoBZOX5B5m7/u1LpAsRGNSS8mPeWAJsMDbNC
TniReOlhRPs3oZ+uW2mRhPTgoFHJO1S6dNX6OvWYQUTeZtz1e1DREZM1b9hFFGQC
TIJGDQAWRZP9HAG5B+QkQXjixdAqcUioMzlo2v678xVv4KEjFBv+cUXl0hx1uwU6
Pcg5rK7M6z+zYI98A7mDw+51eV9sYjQgRF3Kz7ITYaF1nLsvVZqF8yl1/Rmdhs/K
xSVQIqXyAoqqYkO2pd2D3zcZ9Lsu3PrlTIamNHj9E++OSHVCO/1rgqw8Ak9T2mzf
kP+0ZTr1i0fOqUQ0y9nX2h0mqH28mphUkxfb9MhIVsLboKPDEtjg3lMIUDOKgOkn
dBLK0DkL2Wfu/ZnpuS3xPF58BQL3tBvFLTYAH1VKTV2WYfqLFL+A5eiSkBA8Kh3U
wuAprNex26YJJ9CWJmOuWOm6RxESogzkVRzx7RQtCd7w5IfQN3YfiLDLbg/KYnkg
Sz96jqdnMhrHJjrnp29zC7+3lFNjH+w+mszVCGqJ6/CvALYi5KzLsbhzyVvHZnCj
iktavwB0YWYkE3duw0Ju436Uwxsgx0VoUPCIv79fQdan9YdM5k4dnDPWBKIFq+iL
5y5FEe0lfgBkdws+CNSHx2XSJ+OdWGjctv0WcI9QzY1kQIsvIXTcktSoH2FV2vRz
9gkVu3rUp3VU8ZPJbNUjX57sjjToeTHrAFnD+634BFmewD5tnUErgLF5e/jvl5CK
GtPgcGOHhU0th6xjAxugzI4mdZ1KMOiB1+TYH3fxsy8xUX76ShgOMFUyiiMO96za
voHEMtGxrragW/92o5yF1WRr8ZS4g9LR/RANqlFC22rFpmmSVd88jGo9DLNjYxvh
4byb/JGcfiixcjyaTXNWkPqwBmg8wwbNlxQC7sHVWFPZ8YOYTPPe6eqnJUTrOjs3
QWwt+GTw2fNAFCwuHT51dPn0QbpQ/DYVrBQuElifiCoIaEYAaAVDNJ8UzZpWNeNt
+BeXzaMGmNNfHCWJjIHITOPpGEVG/SfnculPlvt8ttMbOOP4fraithBBr52jLhjY
gfdXTIHJN8benswlEAvz+LoAEy2CG0091NcVvi3eWfYbnTSeMKv7SQ3w0wbEXPDg
ibp2fIbA/F0fqTNfXL+k+cIxIVhfHTbk4Pwl6xXx8lwRKKnFK+/Iff6LTn7AJdQf
7fg0rbV/q0jcI9qLOCmsH5u79Y+E9n5wPZfhuiearJE9oYtvSQeTZDl4kMV5AGTh
eYsPV/qVjQhD5GOaejGA5eoYm2zhq+dU36ZtbMX63lFMMYBb3+/Ic8qsBsmuTxk7
xxGN3tZLBIIbHxs1WkBYe9teV6zYjC46Isq8LhxIDW4bI0kHCXPzd5+wE7ph6lxu
Tobs67+1hwxNkSBlh01hU5k/QsqcDkn4bJyPyuSiG4rrQmIeg4aXxd08zVuoRZsW
DxRey2NPW3bAkYkLK5ucEv+WzX82WAwnezVVs2OXOxP+Ajgvl6lmjDddADQ07Ksf
vc3lhejyLMEYBNWnzYd0grXR5XbUynlgW2XlfJQWS0szpoaLo0mYhbv9ecx3be5Y
FH3ugBAXoqzjO5BrwDwVUJ3yS4V6lw5LoGoPfDICzuhXw/N6X58/kuNFcx4DuAE4
rs+gBKq89gCMaDKpT4ItJhehDd/QRKsO/r6PLVaaqeIYpaHkegJ0+rJBGeE/pk0l
qjTwsGHTdzWR+BvfH7AcQOKzr+hkNvT2CPddgQa+KOPBE1H1ZI0q3FG5w/ux92ok
fNVwKJmPl4Ee9LRfxlatCAwMk6lFO5Ox24yth4FTkk4SRy+nbHu88Z3wMP5f7fC+
g4prDjdJu7kq22bjMefQQRt4TI76OMbnZmvdPOSfkkuM1NLI/V3t6ep20XSSPuef
gpRPSH9DZb4+p9dPOWwK2RrgAC8Ow5LgyHOD0GtyJpGpfzZu9TvX+afwt9VmHZZw
wYtrTOEcEiGmlVfF96uTlR5GdyjFY9jdy5zaPNrSI/cLm5VkE8C0MoFhXIwaHs8T
qUY5Bk52Nx4PxlHEe33Ce12shXgxMAiTIaWRSyelHQzDuMZAMibY9CvA5JUHDlFK
oAW3B9JnjP5eCbQaZkBkEpW8PrcVHzpaK7179No9c9gaMC43fdNMJnI5H5IcRIua
ww3arl+P0BJMVQVJd9/pEg6pAEfNYfuzfq2AaHxMqjC4QVQqAsjXKUd8pai3jRgd
uXZnzY02+YcWRX6Du4uesQ==
//pragma protect end_data_block
//pragma protect digest_block
MEYLO5ITOuqlPGfd54pu82vBlO4=
//pragma protect end_digest_block
//pragma protect end_protected
