//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
UpB/1v6M1NSEIZ/jJc1pHhk88S1PEQ0KWMUOefDtW7AWgsO0BPYZ0X5A0t/9nbbR
I4d4z4oD5rrbAAXBu8ezzgM8hRbNz8a85VoOlb0Vxyb4vbNkDgY4qcuoYihlJh+E
3haNH/7qXUhlvb04ZDEMlsXVYkfeG+9jSFpyQHK5uq70b7jUBs1Zd7Qhj9E/jLb2
r0nkp/YYWu4UUhBadrwCEJHTkDoFy40jlW8soi25wnaNW2NbRaT0642cDXUSe3dM
1B2ApnREzVxc4pydlqFIlS7FFZbNeuz1V5EC6uXTztE+zZzGm5p8C6VF5OD7nyq7
Bze5BKh+e+/U5aL2xX5s+A==
//pragma protect end_key_block
//pragma protect digest_block
prgLtvZdIMUq6qjtsW7FS1dWAqg=
//pragma protect end_digest_block
//pragma protect data_block
tusGJSrYZUltvAyg5FRhhtqaxL74+ODJ2qlWJKCawCs5UFpAt2W3sLPmqna2cei9
7dlvIlwKWedM+dSq4pmCDYx/4ady9ipdNagwpmHo6GcTa8SfwdqguzHn/G6uDT6L
ha2bx3m1v/FpNtZImJxgDjfDoBimkqqJuXmWWKiUySpgl188YOcrUGPnhqx+jDmB
LghZO5KP2nwhasf88wHmIfbxbZhPftoLehH71jBrZ9I6vbk0w7Lv4I55Oko0aEVL
WEAnhJH53qWhkkHcAc+um0fXvUQHHVBwaK2/2tM+t+nnKLzO755q9Q34TtsbqEZt
+/vYh6tYMJ5QxVpwpMbXY/PNi3AvCfId7nAy7tEzcC5xJ7U8pGTyuvcFcpNT/piK
vlVbuYmOntTmvuQaoO/jxXe15/yKC/DwTJkwm8iJEXx3iS3U675KETAnTjiNw4aV
AHg5GRyJexHWkpoI9fvMgz6Apt7FZRJvg6sO3NGe2uYPOBlkA8HA4T95ES7gRj6m
+ZJ2GwlCqF5tEwKN0BEZO5MeYXKLRVfa8oRXxTxOxoG/bP5kpRlH8PGGgaK7ENWG
+XOhn/40n+tEUGaEANsxQppadAGxxMF+VdVtNpn/Rhhv6VAVCM99bJkFeilIbFt3
2E3OVN7WuhcRTVjr1UZRs2ZsKohhoXQJpEW8sbBsNShTa7DPeFzoUP+FUqQGD5L8
9BDVHHreow9v2WD9GiFglwolE1NjBOkGcEuOR3tRdRi2obJxzmBdFLBdqZNiU7ZM
vSsH/Zzd3lDEOnROSQX8hQdtwzEPv0E6rllR6fn2kEXSxSBr1bY8SsqPzTPANCS8
kDUTcouES1BxFD6z1yon7JZOa3RhDcdYtiTZj/eYIjBenXZNhJGDo/feMPJgefaD
GblwcbaA0bDR8w4BxEpAazsUbNCP9buw8NIK+ZCZAsup26YShIbI8nPzjZi14NmZ
Q0niBoeoVCyNrQ1ULNIOWZjvgb9TtsRqIjpxgINVZPLPnkoYpXd/iNcKkP+zHNJR
jPRcFKzIDdZOFfBcn0vxMvDfX5rUPi2l9POd1qhBgZE2U9cop6FH1arqa2cpzMEF
xqi6fSEaEJLCnD0c32g71XBTa0yEMsk2T2z23h1OucrXPk4saNMhkTFbPxEJMCE2
oTnfpCVnd+xZl0a064Uj4psBpXvMKFizVP3ug/1zZLq2xm+ieKG5TBmPg+U1JzWx
8KkFs151SffZI39aFQJqpKxVXjQaRvHvqVUaJvo6DQP3nljGjj8gb0BkCtVbLPep
+OK4ussbHNnMNS13S4Lt1Dd+dXR4YEdBBWMnybss47779mCsGnuLgufGg8VVp9nw
f8zHbGhJXMtgvPY5+JxxBjCCWA0FnhYxbelr8q6GiBI49GeoWKCS8eZJxOkxtSwb
Wp6cdu+VJYertxq03itodQgZTt2mO+1rInGSy57xQydKd3nhHFgk8rBhEDHw1D9p
08GIN1UQP6ZV1TN9XQ+xbZ+iK1cDFqIHlVPN0IYE3bL0W31WAQ0w0Hp77c9NdedO
VtXfcjjfQVlBiN+05HptM7PzCPULYG29MDoRSVvcGSHIR1jJ0ZafHxiI2jzeSXHb
ddU0g+5/gfWKrALZ5DnZCi8XWwmU+1UgiqLF0fUWfRZ2VRzYBovy77J3nYKItMSc
fpyDJzw9qF6WtMyHcEewFz6OkwrEs89YPWlmQoZiEnCm7XL8CTiDLKb4+aN/aQuB
GjkEV87wJ2lsiV+18/SIT46q1u/ifmlE/Phe2RfaqBs4NR+z/oSaJJ1fZK7r58Yv
gKSPnY5bD+oWpzfVnZod1pBv1nAXjNqvkdu5tV+72o93HqzGzLCZYO8w/qht7PoL
MlxAVUgQf+079sn5TgORPhsXYSGQpKfUPb4fmICjVuhfZalGX0znjphEhLKJhDLo
UB3BKyOpGNchDz+4GBH6yUDkKSz0aTv4WUxncOMPAO0uDqxlJBRlg1AxPCDgbMOI
jX9lM4t5jcYviiufPx/TtJpighwP/5f8a9lUa01lQrH+hJfp4qv2+TBurHvA/2SQ
NFDXNl8i4VmlztTCNCZRxQPuFrbbFRfBGroTTt+tN7HOU9bRdr/2pS9yjM9wE/uV
wTuK1sR7bM2G4lcngXBBdY1LzeUY85d+9WWNR7zNuNriWkiZbOnc79BDG7Ke3GoC
dIkziz+gheQqsfp3DXtrpe7PrHL5eqpBuuLFu08PIPZu+wBrEWQiuku/Tqg0g/k9
b6Yqrb168DpbDzi0+OoUeoejqZKUdQG7QfnBmuHoAIxr8JGOUNuMfOyUIYZ4YATO
oQ0xMNLvRSxiJfRCEBu5juxn+3q3xME604O2tloy3QxdvkEASZ8+oHPFYImWSuwi
pBxQyDb1/Zn4IMSyQZM++t8M4waylgQQLjrP+pY2W7r9IDE72WuGH3IxPel9fD+Q
Hi1a1XhjpOEMwQJhSVyhKY0CIox+aj42idSi20rsVEBmylh38FQgUyRTLn3gitqp
+W+xRjjlfXHiORWpEYom+KMOczZsIM8SowIJb61dx3sdMDONUS2Nsbny51rL+ziM
9Yub7S3ZyAAr5oY3IQGp6pNbkTYiL77dKun7K0dY4mydR2dQI/aYZXf1JeP2WK2A
MVIHGGMipz+QeWZUHgcCEzcsuvMRupY7K6Pmo2kTNQKpHOytkYUG+OZiEqkNv6IS
kf8IpeiVwXpAv/lWs6kZVbWKWG9zD0FOTVDhlTFFKri3NuZozIqpZmIyeJOA9npZ
QceE6qCbJm4ja4Ow9K+Gs5+4BZyV9oxSQhOhZJ5z0REjbNwhU0Y+veYptBQkupE1
Ynrb6HLW88SbYpRlPg/+6rUdU7l1MFit5846XGLk6XEH1GjP5RF8xt3db6LDH+V8
rje0pzHm2ZUcuBVSD8Czck3lRBSIL1SH06WOjHW6aTSC06i6SpnMzLyhD1A3FLDr
NgqHnIccGcXUTn8wJvzmYVKOtcfAFoY1JufXZT6RFGmwLrT+f7nQ1pzVdVbDgadZ
mwrPevT2swJTOTBK1nFZgIMEcOaMk1DFYUNMrNkIIq+WvSWTqq753Gh1UStUngZu
vypNQT0XlZyzbgw+iDrfDen2zOn1J+h2JtY9uNa9vEjxMX1o+oXBbII/kTwYeevZ
Cic5SjBRNKH3UD9+dXR+GVlLzea65XdFkVHhChzzhc+qPil7Ohi7w9buxKcnJBWm
/atO4rKwgjHuzWHtgo5AJXNi/YBnYwnlMMw0e+h/6EBo12iFFhRnW/PCr44A7F0W
PKq5OoNpboybOBqwHFu4iLkKDFMG8Yfy8avE0q0xURwWAWysQUegiHhqW/nS4B32
yYIFOxagY8epVtKDVYsrQ8n7ecjkECgMhY0MdQw195h3ojxYw9Mg1njxvAPrs5e9
y7XVpSsPUdIQgbeqffDthyas6414iodvX/4fO8oCAm24X0RMxSoiHLszPvmIbzzR
EuMaobBlbY8ZY7/2MoB/U5pKCQLu4UClvPjBvRzJYULsyTnFYvKNHPhy6nr6ZUjW
wHkvqqZNm8tuZ8XkuyPiZiGrLySJ8iDTBc0igd8oFx4NPBe5LU6xbNjKR6gIYNYl
WvEXLO4C3V8e8Lb1ed4K+oDqi2iTUe2nEzNceAUEd8FSTCSiwOCfZPrkdY+cKxwU
2ZbVDpuPSlWaAFqXWye21IDotM2TGeSHkJCIPt+eMKaAaO7yGyFAQx4v3woyk68w
FCRR1HGQKdi7VEoiigwPrUpNsRlsE8l5gFLcknREB9Do3mzWSGS3UAlnm6Rp8Ex4
16swtPZ9xckJURenCBY2aXtGg2tdDc1hJD2WTkBCu0wu8UH+f5rTEQAsJtZ2XnuQ
kvgR/YBGv6kjtvvRZJC2MAsvCuQjl5HMn3RnKae+tCfPhh12Q9UM+m2kzBlqCEFI
4oVHgyJE+UCjHj2QT5nXpEUiD2ZJ6pyu6MNqtrcLbM7I1bVroI129MlYPGCqVhOF
oGE5hvWbscm++C29qZwL6rWv0+W8l9T7i60vN5mMPH3LzghFgrOFQfpridzcXsn1
ePAf55tH8+ps+NOYp/zc9YqEh12il3mnpr+Emz1pNHAaQOUhiNpEe5MHQ1Sq7PkG
mnC4wsDFbSAiLO2UntRZb74Jlg0sAI+MdFCkMgF/BioS7uY3bH90poRRg3UByLFy
PB4Sir2GPFkEwfE+Q3v9TqS+ACtL6iBkTowjlcAIJKdFcVFXBWSJrSHAUr6Pz0G5
cUW0MmlV4udFiCmuYtXij3LvlBWBd05Onz9bn9GrAIVjXZYnkEnJUTNF1Aqr9O7h
RbGpNntFTvpWLB9LCnWxIEFkow0AviOX94LlO3BBwSvaoNqUMp9qGter1BBJHICk
xSq+LPIN0kH+lttamFZUswe65EvUCS1jGW0Lo5kc2r5Xg22k4NurnNrKPqnG6YLy
qeR47X2J22/deVJD0X/xgnGmy9QYypnNKNxAbLFS4g88uAbDV/OeSTuXf/w2xvq2
afIkPcoIybB9vRBXYllJ4zM0QVf60muGB6UJpmDh49JnwxfHGB0O3JMJWohQR3UH
ySFRvsqmwZ1NXBS8Jt3SGguSrX/veZFCThfsHnL/dIs5T7UB8KgTELTc2iWdn9NP
iVRvKLU1goVqm9JeJ/B22lD4ryDTrft1d0H/diNgbPHzib2KaF8H0fQPxbacb0/C
7gRuda+XjOKvybxrA8706vkJNipCclPuuuNxbnyQQYXE5LU/MkPabhvoEQ684IMr
cWtcjfOtFNRr+abRNoCWzLDc65a6ycxWOKcU7xhZOnuy+3PSwpQtvXL6FmX7PMf8
HdJl8RxPdrf1W595bkXubwQYOKzUYiN/Gd13Tvt3jWBcFF6tN6Y+MUfdwLmwnsYS
qiBbkd25mBl5yQXBS5aQkNxMuNgAG2uMmRL/DElGTyiQYzUEjuj4Qmx5XJnT1bzD
Voy4KOfAK1goEb2Bm0QIEyMrwX4hq6rpKM2ZYGcZEjdBdP/ESn1rs5dxAwFQFs54
J19jPFwpUgrlnJBig4l1Bpx5ANcFu5HXfGslyvuIGGa84A62e+OIGxNvlmQZjq5y
kMMP/6MHRnyD34aa/uQQkdd590DpwckQ5HKMzsGdctx6Heqn+zC/H8MYbO6Q9aKG
j0ItmKI3VGWEstgLlFOlstnnqaBGvo0SJ9PBbP97gw+XPldx04RWvMTH1COTMp95
/fL7h81Oh4xW7wGXinRlkycdR68pnCQy0049RriZxRgwURA55UP1y7ZfJ1pge7ri
UFGr4d2aQEOLBU4ZXoGW1Z9WftUiRP7VUSGlkSgSkulguFvlScBvgFUWEyB2wQrv
O57fNiTybTT9a0qxXQTJhz8UtrdTC1P+SzKbheaZKZh+CkmfkZ+G/VLKpFjPtQy+
Xo+B9fcgmV4Qh+zT5SaYXK0QEfrCxIMKyUQtNRZsxM8EY/rhWkYo+fKWmWPzW9Jf
3HzhMlWxKCYWVJFIzBN11mWjyAH2rMEL1HFJR9AMxWW4gQ54lsWLGJKudTEdfb7x
AnrcgFcCGyCLaNiAnQyr50oSAM3ajhMdIBXkd9ogvLMP0z/nTMcpi1Z+k1DsnZE2
1rskF8dMETB2TNlg0TIBsXciDDCc8C6SN4HoQSuuq5jFGBdhVJkIk13y3BNbjUPF
lbhRlZR7NV58SFUNN70GkkSsU66sUF3g1CrcYQsNxX6Cs9g/I9cLnMSw+ImT6S1R
jCbzxVJtcXm/h9VObJrdrB0lSKiivOPkf30KJ4z5EVnGgGya9j9ZBbAb0z9qc3G5
m6rtgpVbmaKgGkQuBsWtqdeUZBbHxOq1n9XA9k5MPVOZBWvhlTHf2mkYODCSePew
IpgZUN3KdlkkGlIFO4/77cKOYXccJNtb5cENpx+b7hvec3ezeSDjUVrs0drZRXA1
e4oYVKkSJS2IqMQOp8fxVbbuW1bl4S+rwfxbYu/ZZoHxjJgAYAC5r/0rRONyzSEu
3tnBmQzrtdSblfQVWv1WqFPFJ4JnVFJ9OOisOmXR+m14RBUtCwkkrOaIm6Auf77G
0IIqCU1ZICXtgqdftR7upIr7/GfFIrk6W73Uv0IQP/BnRWZ7fmaZuOiIlqugkpUB
w8CJ5IG21UAPdVkaU1afztga2GdKO4PmTQHVuiKC3K01Q6bZksNgdLvMW5+c7gcB
ly8SsUqEAO4mGjJxKF26fYSK51IU1sTSABRqBGgae2LtC6UIxS88ETG9f/Z3DaMO
Ah/w8KX3kR91rAbJB3DJ1H74dsPdyUHAdm7m8sOfsipShjU08u6yJqJkSUmthioQ
TUTftDYO5rl8EMDTCsBXi8zigoSpBBlLCK/F9pu4R/9VGFIGQF0NADifMqWoXxZj
pXJU69UY769wsHwgZQQ+qzNQHDa0EjC6z9uwvc7gnI4Xp8834TSNdByxfLk7Estu
8Ikc2CncRvVg2cV2pqwvWKz11NT50yzGNFgrRqyzAv7OtbTVs05z7k/lA4wXbJqR
l/0dr95wckliplgQDlHaQZ/a4zm1mRZZimOP6A6rwcDYegf/3rr5AF6/9EpPamux
bYYaZqAMkNo/v7IwWbchFWCuzOhXGRQHfLXeykal2ZnrB10KdwcvB61yyQoWyaQ8
QEN8cYfH36KHYS4V8oymCytV+6JOrQuRwIBD5/nRon7R6ZolHTI6z6c0wVJDqw1c
48oJOw5NqKTc+5cvgjDkEVF5kwFutRKVL3qcf6qZMeSMfVC/8VqTLXnWBhtJiyrI
vrczSjmCzRUAxjqHYZtQ0SL7nlf1OPZuXykHpRJF9jPg0V8xXVFwlXFTa5h46Y00
a0G6rBavYw2bbtNnFFWAxFrnpxdbWeEuvDzH8h8/S4m5YO1YHuDRw4jZN/dcIZyj
AothXSaWnEJRT8AxYiUed9+3CYTBlgjkmjPhDO/8pAILmfH9UsqRdR5EMHP5RW4y
ZuTwyit9a7Uv70CewUhFrQ8A6JmIkF5fylvrH5j5Z6wIMN5AZSuhqZNSYmNQ9++U
m08rDD4To3XttKdR266MNkyKaevgPUGAkesSOhb/oXkBTr2IjpJGtSiBH1eh0veE
Y/ya3Ye9wu2w7U5wGAMkYTHbJcm97nFcWujqWMB+DaKec7XNM2xzNABI9BY1OcD7
WOhLKt/9+7jx9yYrHLB/XSQiF6olaOM51gfPwE8UkulEIEBELO1UQuf7TcISWvdv
KytCJZ1uGrvPRm6Y+RqRGyVAN3MJL3osA4Lit0rO/BTc7nQkzbH4DhA/ADHFsF1X
bA5v7zVWEDEBSG/jfaBvnPJy5E35RCaJfrBNcAHNof453+ypKucAq4RsduomE43P
M60LnntkygmZnvfgTJOPcQ==
//pragma protect end_data_block
//pragma protect digest_block
TJIMeqJ50AvuMv629UyxYHuB/dU=
//pragma protect end_digest_block
//pragma protect end_protected
